<map id="enemy_movedown" name="enemy_movedown">
<area shape="rect" id="node2" href="$group__xpm.html#ga8b990eb150243edd20fb9c4182748528" title="buffer_destructor" alt="" coords="181,5,300,32"/>
<area shape="rect" id="node5" href="$group__game.html#gab806d0bb50ec52aaa6ad9a71a2d3a05f" title="Says if there&#39;s an enemy going under the ship. " alt="" coords="209,56,272,83"/>
<area shape="rect" id="node6" href="$group__xpm.html#gab41dd197773f68e69e18c73a8119ba5e" title="object_creator" alt="" coords="189,107,293,133"/>
<area shape="rect" id="node3" href="$group__video__gr.html#ga1cd7727ad0fc3fe3ffbbb98cd9115c1c" title="Returns a pointer to Buffer. " alt="" coords="351,56,424,83"/>
<area shape="rect" id="node4" href="$group__video__gr.html#gaa55320d571dc2cb8179422a9d8114de0" title="Returns horizontal resolution. " alt="" coords="475,107,547,133"/>
<area shape="rect" id="node7" href="$group__xpm.html#ga05b2c5e4dbcaffa701703b50a2111783" title="read_xpm" alt="" coords="348,157,427,184"/>
<area shape="rect" id="node8" href="$group__video__gr.html#ga36218c155eade74951ce7ffd60711a9e" title="Returns vertical resolution. " alt="" coords="475,157,547,184"/>
</map>
