<map id="start_game" name="start_game">
<area shape="rect" id="node2" href="$group__xpm.html#gac0e395e7e8c65b90f0680c7a917f1acc" title="title_creator" alt="" coords="627,347,718,373"/>
<area shape="rect" id="node4" href="$group__video__gr.html#gaa55320d571dc2cb8179422a9d8114de0" title="Returns horizontal resolution. " alt="" coords="988,296,1060,323"/>
<area shape="rect" id="node7" href="$group__video__gr.html#gafa847549e9dc6e4f49f651623bc456dc" title="Clears the buffer. " alt="" coords="806,448,894,475"/>
<area shape="rect" id="node9" href="$group__game.html#gaff72f275b5af37960b3baee51f855041" title="Makes a game round, where updating action on screen. " alt="" coords="177,397,231,424"/>
<area shape="rect" id="node12" href="$group__xpm.html#ga8b990eb150243edd20fb9c4182748528" title="buffer_destructor" alt="" coords="613,195,732,221"/>
<area shape="rect" id="node15" href="$group__xpm.html#gab41dd197773f68e69e18c73a8119ba5e" title="object_creator" alt="" coords="316,245,420,272"/>
<area shape="rect" id="node17" href="$group__game.html#ga425ea598437d36368c0e136f2be75a61" title="Makes enemies down movement. " alt="" coords="140,201,268,228"/>
<area shape="rect" id="node19" href="$group__keyboard.html#ga6d2cc119f3d1b28fd79e7acf2f4d4596" title="Reads scancodes via KBD interrupts. " alt="" coords="165,600,243,627"/>
<area shape="rect" id="node20" href="$group__mouse.html#gad34fbf075c41898c2120ed2d0ee6b20f" title="Reads packets from mouse. " alt="" coords="156,651,252,677"/>
<area shape="rect" id="node21" href="$group__mouse.html#gaab4aa4fb914d5e1046d1391b97091546" title="Checks if the given byte is a mouse byte. " alt="" coords="149,701,259,728"/>
<area shape="rect" id="node22" href="$group__utilities.html#ga88386f4f23c71aba0d4e995a5246f981" title="Converts a number to its twos complement. " alt="" coords="141,752,267,779"/>
<area shape="rect" id="node23" href="$group__game.html#ga1fd9e64dab3abe9facfb4dd7e1267bae" title="Creates the pong and switches game state. " alt="" coords="167,340,241,367"/>
<area shape="rect" id="node3" href="$group__video__gr.html#ga1cd7727ad0fc3fe3ffbbb98cd9115c1c" title="Returns a pointer to Buffer. " alt="" coords="813,245,887,272"/>
<area shape="rect" id="node5" href="$group__xpm.html#ga05b2c5e4dbcaffa701703b50a2111783" title="read_xpm" alt="" coords="811,347,889,373"/>
<area shape="rect" id="node6" href="$group__video__gr.html#ga36218c155eade74951ce7ffd60711a9e" title="Returns vertical resolution. " alt="" coords="988,397,1060,424"/>
<area shape="rect" id="node8" href="$group__video__gr.html#ga5c30cdd3eab0edd2734ab3871f7000c7" title="Returns number of bits per pixel. " alt="" coords="968,448,1080,475"/>
<area shape="rect" id="node10" href="$group__print.html#ga1243268c621c2049a41956ccfc934fd5" title="print_info" alt="" coords="331,448,405,475"/>
<area shape="rect" id="node13" href="$group__video__gr.html#gabdd05df698103c4641478f491e11e284" title="Copies buffer to video_mem. " alt="" coords="780,397,920,424"/>
<area shape="rect" id="node14" href="$group__game.html#ga9a691a2142903ae9009a88a62464ddd9" title="Says if there are still enemies. " alt="" coords="322,397,414,424"/>
<area shape="rect" id="node16" href="$group__game.html#ga8aead8655bcc62fb760afdf2fe161ab0" title="Destroys the enemy hit by the pong and desactivates it. " alt="" coords="477,347,556,373"/>
<area shape="rect" id="node11" href="$group__print.html#ga4316256507429b01e848fd72e5fdca73" title="print_number" alt="" coords="468,397,565,424"/>
<area shape="rect" id="node18" href="$group__game.html#gab806d0bb50ec52aaa6ad9a71a2d3a05f" title="Says if there&#39;s an enemy going under the ship. " alt="" coords="337,195,399,221"/>
</map>
