<map id="is_enemy" name="is_enemy">
<area shape="rect" id="node2" href="$group__xpm.html#ga8b990eb150243edd20fb9c4182748528" title="buffer_destructor" alt="" coords="132,31,251,57"/>
<area shape="rect" id="node3" href="$group__video__gr.html#ga1cd7727ad0fc3fe3ffbbb98cd9115c1c" title="Returns a pointer to Buffer. " alt="" coords="299,5,372,32"/>
<area shape="rect" id="node4" href="$group__video__gr.html#gaa55320d571dc2cb8179422a9d8114de0" title="Returns horizontal resolution. " alt="" coords="299,56,371,83"/>
</map>
