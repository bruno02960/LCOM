�PNG

   IHDR     =   �Oe^   bKGD � � �����  cIDATx���{T�u���ܸ(r	��H��
/�f����m�%�~�Y��R���n��L��w�l�mw��JWL��RKrI%n���"?T@P��3���g`��g���N�3�7�|���~��B�$	DDDDD�k(E """""�b@DDDD�˰ """"�eԢ9���55hmmCss+t:���׷��W(@`�?|}5@XX���DI����z46��ܬGc�MM�0M
�F�B@���q���D�%�"���d�d�PZZ����8{����p�b���v}�F�Bhh ""��#"�{���!aN���w��%de����2Μ��ٳոq�ժi��44(��; ����qC0rdT*��A�)xw ""��������(,<���r44�臡C�#::QQ!�����w��@���ѧ�/���������>>�G0%46���j��+M���Gmmjjp�\JJ�p�BL&	�ၘ4)S�ǔ)�1hP���A^('��w���S�����q��������~����AP�?���J�DccZ[�hnn�����p���Wq��%�痣�����5k,�����1P(��\�DD$g�T!#����8�Æ����1?~�0��"�T�n0��p�l5�����gq�X�뛑�0?��HJz !!}]�>y?I�p��)l�|���HH���G!1q$��#��Fyy-��;����8Q�ѣ���<O<1�� ub@DD���;��Ev�������� F�pΠ�^F�	99e�js�o_t�6,X0	K�<��� ����\�x�����G�!1�^,]����!.m���"��������8q(6mz�G� � ""���o���Ą	C�b�L�+˽�:����ؼ� ����+�`Ŋ����uԳ���r�DF��c̘�nm���"�-K��uش�9<��X��O��"��������vm�ǪUO����EG���`�֭G��?�ETT>��y���d,=� K�n�/9k�̂�����`0b��L��������ܹ�� y`@DDn%I֬Iǖ-�a��'�xq"�jϻ�IE�U,[��'*�e�+x��a�#�8p/��	V�|�?.: �����/l۶?':	�"����jݺ���#���1m�H�qb4��b�����o_�	���D2RWׄ�S��s�MĚ5�Dǹ��o��?�AV�*����� ""r���,[��-[^�#��#:�SH���+Sq�p	\��@ёH&������X�F%:�m�F��>Ę1�x��gE�!<��+y��Wo��7�������#�@�o�Ng�a
�7�AA}��[���L�9S���\�[��FI���f��J�Ě5���EE�U�qH DD�|}��"1q$�~��qqo����
��=�;rp��u�qH23��w�Õ+�x����o�\t��L�8��"--Ot��5#""��~���g��fČ��yj�$�gϨ�&M���Ñ�r+V��0���)ÿ�}[�|��z�.M�Jվ�U��O�>
��#9y��(�f,���%#:�6_}UI��q��` ����t>�#GJE� 7��k�ܹAY��th4��>.I@[[����/2�Y#GF���&��ҧq��� ""�khh��� j��s�U�@�[�Ņ#==_tr���+p�ԥ�ז�uHH_wE����!0��r��ၢ���y�>}|�_4k� �F�
&����D���O���?��t9ފ���ܽi9�v,�����j%���Dhh@������mnL�zMM�^w�Ygժ�����bW�U���T=������>����� ""����֭�@�Rv�m�JN�Lt�S�.">>Rt@�Q����b_W*
��3$�˯�_??��ȯ@!�b@DD.3v�@|���1�B�$>|S�z�C��v��X���f/�U( �#EE�3&�b�BދE �ԬY�a��',�y����͉\#+�����9s��($Я�ƍ���	�F�$�#�~[��.:	�"���\.9y:f��Zu�{&�$ ��}��A$%=����QH �R�?��yh4*ܺs�h4"(H^G
/����<��($ � ""r9�B�>x��fO���"7���x�㢣�DG�`��_@�~�$	�ב���-��7C����B� ""�����������>��A���E`*�UW�������E�"..Bt��ٳ���'G�v�P9	8{���?`ɒD�QHDD�6���ز��no�IZZ�X��DDⷿ}Rt���ߟ��@�΋n�tM��of >~ f�%:
	�ka""���7�7�x� ��3oj4���l���u�䓅��Q��D2��7?Ij��E.E@jj..�ƍ��@��B��7UUU!99F#�g���XlذAt���v=��y�0k�,�1쒙���[���!ԙ3���鋄�*��˳�u�`P��8���Я�^taT*6mڄ��<j���(--uiǏߍ�FL�|rsWT����С�.m��?�0����HII���裏�3����� t������={��(^I��`�p�V����c۶m���e��HII��u'�N??�}j�$A�:��Z-�mۆ��狎b��=�\%I�^__�����O>,m/-�|��7]�L�2�ׯ�a����#x������c������EQo8�ē����O>,}�&�������a@DDDD�˰ """"�eX�2�*{�1��wE���p�Y���}µz�����e^���F���D�pW�Z��[�;k�.z�o2I��)Ò%�p��E�Y���[�q�ؽ��
�X�����bko��>�׷a߾X��344���=Ѭ��<��55�"--���mm���8kq9�Myy-֮ݍ;�E(w�V��7t��'/"=� Zm.�\i �Ņc��(��H�ʮt��� �Z�N�Gp2�f4�p�H)v���_Gss��f����{�#�=��6|��i��U���O@�o ���?ETT��t$Ruu=���Zm.���w���ܹ'�~N+:��:t�=�:t�{������ki����k���5��=��5�����v���k�Ѩa0�?(��O푕�B��c�������tl����Ξ���u$[O���{w!RSsq��%h4*�F�Z��}}�֖;u�w�~��u����ص+׮5�6o=����\67���ϱg9������27]O9mmǖ�HO9�5O�{mn���s��h�ѣ�sg>23@KK+T*��<{Y�r���f��[�6�_�R��ǣB11aNk˝\�<w�=9�)E���jsusts�}{���uOm��]{u�ho|t ��������+��=[�Vׯ7�_�:�6��巭��a�jNw�0�'�QRR������ҥ�]�=��Os��3�����8��9�R�SN[�p֠�Y�Ԟ���^@zz>v���ի7n[=� ����v:���c��<:T���-�I���7p��������co�g8R(�2��{��J_l�~�lE�M���[w{<:~����yϑߵ�B�AFF�����%��xI�`4zϊ��nTT�裯�cG.JK��v�+{����sE�3>�Y,m �i�ֽm�rd���u�+>���ﾻZm..^����"�Ck)o����{����v�^oc�w#r\��-���ו <�7X�|G�Ϭ�h%	ذ�l���+����_%���lx�n�]9���$���W��<������g��ݶ���ƈ�`VC���w����!k/��wWŲZhhƌ�å�5��k{���u�����o8�{�@q�Ϭ]Ǐ_�P��<Ct��\��������Y���ԩK0 �U���P���\��,��<�^n4���[L����*�T*�>���3	�1c�RZv��wظQh �ً�C��|�B\��Ӧ����0���~X�?&O�y�&�ݶ3dgg���k�f�$ ����f��Aii�j��5^��q������_�(�}wu4�է5x��֕��+���ƅ��JBe�U�����[w��ƍ��]w�u�}G=�� ^���D._㩧V���--�T
���U�f�!�e���x�]��>���v���E�5����(p��w�q�{����	{�"--ǏW@�R�h��.�
�Y����G���l���?�:�����:�w��9--%ؽ{)tػ�8��<�䜻yH�|� �A�Be�?L�B3X�TJ��k¶mo�ܹdd 55W{�x�������m\<u�멹���ו&�������q�D%��󑖖�������bĈH��s6����i<�?�;�^�v-Fkk���v�����'o����1�U`��,��{N[uD�)E@�;�t�k���� �_����v�U�EXX ^z�a���è���y�bii��ܝ�Y��]Au7����҆��0o�D̛755���,�V����Jh4�Jܦ8�#�a��c��X�|������ɦ#���>�����Z�i��^�����a�3]Ŗ����9�w��ѣ��f�ϐ�S���dd���j��e�S�y\m���̙c0s�44���'����#G�B�h?���*Gt�C}$��A�������������i���%�X�$����A._n�k�N�����_�{m�E{��p�=gf�N����p�T,\8���u�eeW:Ɩ���u��kK�9s�;c������p��9��`��Bܸ��R��Ҭ��|��k�kG��7[O������y���T*0i�0L�4���YY���]���b��m�$���8�C��aΜ�3g<jk����~GŎ3(��L��S�4�Y�o�'{��0bD$~������{df.Ë/N DG�%8�����x��i��^���^�E� �Ɔ���Jz(�7'O�ǧ���'�h�g��P��z�F�i�F�/y'O��G��	�o8(8��_�j
��MƱck�r�P*5�Ru�����P(��0		���[ψ�#{���=H���@|� �^�S�Q�J� dڴ���Ț��9wgsV{r��"��������O�/:�l��>s��n9��޼�#����	9/s�����<O�>�y9$��Ӂ������s� """"�eX�2,�����z�gee�1������jEG�J�2_��wh�Z̞=[t�h�Z$%%��A��i�Zh4�1�����������" 66 �v�Zק�>>>�#ح���3g��$ދ��ubbbDG�[LL�l�-�-:����������p�'涗
���"""""�UxM Q/�"�������a@DDDD�˰ """"�e��fa��\    IEND�B`�