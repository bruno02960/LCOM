<map id="getSec" name="getSec">
<area shape="rect" id="node2" href="$group__file__handler.html#ga90d3bc0149cb0d2782d63aa42cf3fa86" title="write_score" alt="" coords="116,29,204,56"/>
<area shape="rect" id="node3" href="$group__game.html#ga02fd73d861ef2e4aabb38c0c9ff82947" title="Makes game initialization. " alt="" coords="252,29,291,56"/>
<area shape="rect" id="node4" href="$group__print.html#ga92978930f74831bae9a6d6f22d089615" title="print_menu_kbd_or_mouse" alt="" coords="339,29,517,56"/>
<area shape="rect" id="node5" href="$group__print.html#gae91d4cbee2dab64187187499dd0eecd4" title="print_menu" alt="" coords="565,29,652,56"/>
<area shape="rect" id="node6" href="$group__spaceinvaders.html#ga3c04138a5bfe5d72780bb7e82a18e627" title="main" alt="" coords="700,29,751,56"/>
</map>
