<map id="title_creator" name="title_creator">
<area shape="rect" id="node2" href="$group__game.html#ga671b58f5509a3a9fa692bacccfc32cc9" title="Receives drivers interruptions. " alt="" coords="603,144,690,171"/>
<area shape="rect" id="node4" href="$group__print.html#ga92978930f74831bae9a6d6f22d089615" title="print_menu_kbd_or_mouse" alt="" coords="835,208,1013,235"/>
<area shape="rect" id="node5" href="$group__print.html#gae91d4cbee2dab64187187499dd0eecd4" title="print_menu" alt="" coords="1061,208,1148,235"/>
<area shape="rect" id="node7" href="$group__print.html#gabbb46faef7390f85ad76868944abcf20" title="print_score" alt="" coords="289,195,376,221"/>
<area shape="rect" id="node8" href="$group__print.html#ga5f04c1438b5689bedddc17eb0dd9d060" title="print_message" alt="" coords="593,68,700,95"/>
<area shape="rect" id="node9" href="$group__print.html#ga4316256507429b01e848fd72e5fdca73" title="print_number" alt="" coords="144,144,241,171"/>
<area shape="rect" id="node12" href="$group__print.html#ga2eb771fa3527f72e821a14e413498d1d" title="print_instructions" alt="" coords="424,296,545,323"/>
<area shape="rect" id="node3" href="$group__game.html#ga02fd73d861ef2e4aabb38c0c9ff82947" title="Makes game initialization. " alt="" coords="748,169,787,196"/>
<area shape="rect" id="node6" href="$group__spaceinvaders.html#ga3c04138a5bfe5d72780bb7e82a18e627" title="main" alt="" coords="1196,208,1247,235"/>
<area shape="rect" id="node10" href="$group__print.html#ga1243268c621c2049a41956ccfc934fd5" title="print_info" alt="" coords="295,144,370,171"/>
<area shape="rect" id="node11" href="$group__game.html#gaff72f275b5af37960b3baee51f855041" title="Makes a game round, where updating action on screen. " alt="" coords="457,144,512,171"/>
</map>
