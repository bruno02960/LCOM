�PNG

   IHDR  �   =    x�:   bKGD � � �����  3IDATx���ype��o�r@���+�59DN���]@dr�d}U�u_�(��UkY(]t�"�����B3���E H$� �#�$&��k����!3����~�,����oz���M��OK&��"""""�4���}X�y(�DDDDDJ%: ��hBYY��u�����`BMM=��m�$I� �A�Q�k� t��Z)8=�y�n��ƍۨ��GMMjkQW׈��P��Gpp z�����X�v,扈�m�ʪq��e�>}���r�&�^��k�*���z���D�n����b��_��hx�#�)/�����ͽ���p�|	�ʪ��W�R�G���wèQ�0rd?��;vpqj�tG�!""W))���{�y	99�QTT�J�_��~����{߇^�:�w���ի3��T�B!�S�P*�
��`DMM= ���z����(/����PQQ���
�?_���KP_�����F�Ä	��0!Ç�A����6׮UB��ľ}g��[�����x�����Νѱc�! @�� ���a0q�Vn޼���(.��K�ʑ�y	.�B�R��DT�<��hD��$?�X��SUV�bϞ�HI���c		��1�}1jT8z��K��ф��
���ȑ��ȸ���r��cΜ�x��Q8��˖O�����7�GRR6�v�'�xS����N��UYY�C��a��8p ��~x�������l=݉�<9Gyy6mڇO?=�Z���BT�L��_x����r$%ec׮,�c�����t����\�yt:6n܋�� �û⥗~�9sF���WV��_�:��?��
o�53fu��ȣ��'""���6�����#(�˗O�cС�Zt�6=Z������q'��ƍ��Et,� ���x��m��ǟ�z�S���֮[UUuX����?��ߍÆs�T�Y�b���엗w�ç����K/��M�m�ڱcx�$U`͚(,\8Vt$��+Wn⩧6�G�`l��;���UX�}��`ٲ�0![�<+��/��<������[1zt8���t��It$�56�qc>�� �.�5���ߊ�D2TQQ��3�C���"���_�z�T1bb�`��aذa��8$�2�6CDD6�ȸ�E����`���{d! �
���$�ly~xo��_ёH�^}u��5ض�Y� 0thl����!55Wt��<٤��
K�~���1x��9^�gwƌ�������Сs�㐌8����<��E�S'y�"3rd_���o�f�n44�E�!A<LDDn��k���kg ���'r�)Sa��X��?��m�d��7�`��G0th ���f��d�$(�
l�~Dt��<Y-/�
���êU�c��#7n�
�EGs�+�A�$�����($�ϗ ?�źu�x䑵�������B�Vb��Q��?&:
	��\�U#��sйs ~��m0�L0��P(+�:����T
�ƎŶm�aѢ��� /����|h��!IV�N�Z��N�ԕ���Ap»M�6qq_���
���aV}�y""�(?�:>��{$$Gee=T*�zyu5p�q�"��;i��jt��Qtr��kwc����Р�J���hB�ͅ< ���ئA�zB��p��5�>��<�����}��@�V��n������ \�P�bއ�&|�az�c��h��!!nHd=�Z�n�:�����($ ���Y]�h��?o*�U���46z��D�S($�ٳJe�wt�ۙy���z�/fd�y""2��w`֬�P�|�pQ]] 
����mĈ�x��i�[�$�_�[]]#�f}��읉��f�$!..��l9cݖ�:��1?�:T*���!:
	���S1p`��]nc�M��޼Y���>��<Y���֭�`�����Ş��o�aذ��,����j%�������:ɯ�ͩSW`2�0dHo�QH �DDԮ=B��g/@�T���@��_�{��됒����ᢣ�@��/y�Ͷݹs��D�}��9�]���B��'""�<�p��~�=�+jj��.����`4�=Ft������t�i�(\.L&���f��P_�b����6s�0�Z��=g,�o��JKoa��4,^<	�qH0I��iS,:tPC�s��R)e7,eZ�i����#DG!AX��MV���3n�F�#{��W>G�t�EG!��;�̇����
IV�R�L&��nf���0^��X��M$I�{�-l��d2��ڳ��l޼����~~��"�b֬�5k�j%�������=Ν+��U���B��'""���k��'K ����sG�IJ�Ɔ_bݺ9><Lt���ޚ��� Y󥥷�vm*�,������@��d���cII	V�\	����"�T*���P�Q���k���ŋ�cx-�׉������Eǰ���/�T]��ɓ�ЫW5�ëDǱ���!�h����3�;�3�<��3g��a���T|��g.]ƭ[~���n�[�Z�.�UUc��r(���f��?�0s�\vO1���X<��cn'���رcbbbDG�Ks��y��	N❴Z-ۇh�Z M�>=Q��Rn���P*M.-(\�d��1�}�V�ELLv��!:�]bcc��m��A	��I�̶n�����r�َ��W�va$�IOO�a���ɝ7\�'���\{������ۡ'�3�����}扈���<�y"""""�b������C��'""""�P�*�'O�l���^K����u����&\��֯��זu�k�\�m�l��6#��o� 7W��~����.�d���|��wx�$�9���ᐸc����}t�֥��bk���&N�,ƪU;��q�-���ρ�#���h�ѣx��x�9sUt��h���z$$dbŊx������9�2�Ym������!11�a04}P�����䠪�{��BBB&��� FcS�x�ϼ	���!%%		�(.��iG�裑����ӧ�"99Zm�˫ ���1xp/��H��=��?���l|���tM7����@�^���~N+�Ϝ<x�'O�����g՛�o~��k����|��ښ�̳���z8����l��w:����B�I�t�ն[���|�l�Fji>{����H�������7g�������a46��hn�-˝Z��;?ws��|��~��w�B��D~�5�TJ��M�J��NY��Y�>�j�m�g�o�}����M3��Zm��^N[�c�~����Z���5_{�u��OHJʁV����
��ʖbM�V:uY��m�1�����={N��N�R�^��g�]�=[����)�|���ܴ;�U�;3�#�k0q��E$&� 55uuP*)$<�f�vik�o� g���|�N������8|�<����嗧P_�;0K,�O��6a���Z��sZm&��
�T*Z�k����m�m�gϺo�n[y��e��o/��}�U�8k�ړ�[i�-�����]Y8s��]|�ހۢmL&rr�������lTV�B�V@�k�O{G���ٕ��ӻٴ>���{�R�;�K���5�󟓑���7nߵ��B�����B�j�`)�=�y��
k���HN�Fee=�j��v`渲H�))9ص+�����شLo���do;w���֗1g����;�Y��;�~9ʑ}�����x�^���c�j����B(R˯��T�߉ۢuJJ���[_B����땭��y߉,k?�uI3������g�������oy�ڝWϞ+]��zCEG�� �������;>�͛��zN�k?kc�^�#$d��m2���З�t�g6ϻkW�m���l#I~�#���
c�.�S���tt����Ç?oy�������o_a��=-�q�c��2�\KԶ��� �y�4��-�Y[���E�����H�,��G��F]�;vJK(/���[g{�ly����7{�V��rF�U?:��uu���#Sp�z#nެ��}�T
|��3-��~�	 �s�&I@ee�L�_���ś%c�>���G�:�E��_uB3���_�\�U�SY�W:��T*x�;©S�P($&����'�ԩ�Z��6m�$t�� j{hh���#���Ā�Wo�Tm�0���№��>�t]�;9���f�xk��8�O}{�*<�|$���ر$'�`����i�J���s�̙�ܒ���M�oݥ�Y}�����Y�u�����X�(D�ȑ�HJ�Fj�ɟ��P��/�P(d�>t��̪��_|�UUu��O!!!Ǐ�\La��ݻ��u[]}��?1{j�꩹��;��aa�رc%�ʪ��z�ve�ԩ�P*0f����C�o�;w6�5���iw�6�pa8bbb��[���$&f�ƍ���#���)S	�����^"��;��o=�L��k�ͦ�;vk(Ə����X��i������l���A�3@�$�7�Nm}hf�N��|�N�e�R*�8�?&N쏷ߞ�u#9ʑL�N������1(-�Bjj�H6yyW�����&����ڮY���^���.���t[�k�����q���x�$,^<	EEHI9������ǟl:+�	�-�fذ0�ի��ѣ?��:�۷-���V�ۏǟ��T�����y[������B�Vb����:u0jk��ק�H-]<U{xXzl��i��pt�3�Y�Ѩ0}�C�>��V� h����`Dmm�ӗ��>ksӜ���w�%K&aɒI�|��e\�K�~)&��=�{�5�Ԟ��������������9{�#b��j�#�º`��)X�|
��!%���L����ۢ�
	&D`l��t�311_}uz�&���/9r����6�N��[h5QQ#PYY�/�<�M��i�i��� ?̝;
s�BEERSO".�+Y\�����+�aŊi8{���s����]t4"�2p`O���:YY�HI��֭���>��H �F�iӆ`ڴ!�}�_}}t��E�'8��M�co���q��':��Y*f=���5�t	�s�M�s�M�������?):�l�y�sw6g-O��TI�0zt8F�Ǜo>-:�l�b�	����#0{��Q|�[�ِ�����\�M�y�sw6g-O������"y�� DDDDDd�DDDDD��<��b1ODDDD��^ ������Z�j�Zt�)9��V+:�Sx��A�K��b޼y�c8D��"**Jt�!9�le�8sO1 X�f���T���4RRR���":��b�p�F#:�ݚ�����'!r\xx��v�N���"<�Ƀ��d��IDDDDD�h��y(�DDDDD��<��b1ODDDD��<&����    IEND�B`�