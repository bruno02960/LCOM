�PNG

   IHDR  3  9   ��~�   bKGD � � �����    IDATx���w\U����eoADA�nŭ��ȍ9+���/-�~?[ZYi�f*���Z�����b	*�2D@����Ji@�^��|<x��x/���wI
�AAA��e���+AAA�
fAAA��D�AA�NaFAA�:IC���<w��e��d2e�R'����6L�e� B�% 4`�������;V٥�9;w�DSSS�Aj�T*'==���\����. ;����rr
˿����SZZv�*7��\�B� 7�##��}jkk���	����F��06֥Q#=5���D���z4ib���	�J���YD��;v(��:���W�%�POܻ�K||�ne���IZZ��٤�fs�n6ii���e+i�cc=������1�� �����~Y����@&�#��������?/������
�s�~y8z�ngd����1͚5���++ll���{{s45�k��&�3� � 5.7���ػ���%>>�������QWW���,-�i�ڂ޽[cii���VV�4ibX�A�Pp�^.���$'g���ERR&���\�x���{�����N˖f�i�GGKڴ����[�&�Z����0#� �PMJKeܸq���������˵k)ܹs�D��McZ�4�ή	]��agW�}��*ٲ!�H��0��N�Z��q�BAbb&׮�{�������A��H155�S'[�t��K;ڷo���8���x5	� � T�\� ..�K�nq���\�MDD%%RLL�qv����
//�hӦi�w�0���4��ӥ�~�TNl�]Ν�',,�-[N�����Ҡm[�t��O�6��a��!N�;D�AA����BΝ��ܹ8._�͕+w��-��D���m�۷��{Ҷ�F�.W�44�pv���يi�z���͹s�\����㱬_==-z�v`�@gp�¢��+�f�P(|��>�5k���n5�a �HP(5�AUq�n6g��q�\<g��$&&uu5ڶ��sg[|}�Ӯ��RA�6�=Æ���MHH4!!Q���Y�h..V�°a�qr�Tr�B] Q��A��rr�pt\���v�l1����Ʀ�S�۶m���"�T���̶nݪ�JA�.���s��u���ԩ$$����E�N�����ݽ;6GWWK٥�;��2N��Ahh4ܾ����c�tf�莢�Fx��"�B=PR"��vQ�m���ՑJe89Y1jTG�m����"�T�3�P�K9>�c�b9v,���D��4�ڵ%}�8н�=nn���PSv��B�����{�^&'���=[3zt'�iW��	/D�A�/��>���`��T*��ނ�#�Zl-�f�f&�Hʿ��~�����?|��}Vv�'��I?Ce��0#uӝ;�tm��ԩ����bM�>m��ǁ�][��-z᫊�)�_�?.���/�ԉ�3�ЦMSe�'(�3�P_<-�<NC��ŦysS���С�H��>�?O��
��ݓ�HE���Su��3�P7�drΟ�/�q�Z
��ӯ�#^^.���SSe�)T@NN!�u?�c�ťѻ����G��$�߁P�0#� '����<����-"7����b��˾��������՚˿/((����L^�c��] '�x����PP�}<o���سnW�gaFTWaa	G��p��UBB���*��ي���t�C�����cu�B����kl�x�c�b��k�̙}7����Z# ��TNFF.w��p�^w�fs�^y���q�~���<23(-��k����kch����.���k?r����,]�'EE�g�Uv�J����!C�aa�ϲe��PT<UG7�n���i}��vϺ- ���EGq��UBC�)-�ҽ�=�����++ce�(Ԁ��Sٴ��q--^݃3z�P�p�0#�%�+�w/�;w����,RR�HK�%--��﷖���h�Āƍ�����>��}��`d����.zzڕ^D��q	99EO|�aײv�l������02ҩ�13}����hK�3�����q��U�����בH�o_Gn�����)�D��de�i�16l8���o�9�)Sz��%�?�ss��� <A~~1		��ť�N||ZyxIN�*oI��T�i�FX[�Ь�	M��0��܈�M����Y[[�;�<0M�2~|WƏ�y���֜���j��"AF�)**%00�={.���//��v��;���(cc=�~ۇ3z�fM0˗����`�'�ǻ���1f�K&�s��}��S�y�ރ�R�u�^.P6��Mclm�`ooN߾mʃ��Mc�͍T��uZZY�jjj���&Nt�g��560򟳇=����	�P����8r��w_$00��)��9�j�D��\D�"�\������#�5��W��{�n�a>�x��;)�<��0#�{r��۷3���KLL�Wl�]�_O��X����f����������;�&4onZ��^�ұc"#����Q���j���EZF�����N�u��v�8�޽���,�[��|��Hn����B&<��E#V�Ü9|��~&O��С���ÑXZ��S��3B�RZ*#&�.��wO$<<���
K�H$4o�������k������������߿@�%� ����lv��Ν爎N�ukf��ǘ1��*�B�5on�?LeҤn,Y�}�|ƢE��1���zVO�0#�Y��2""��CKxx"��ɔ��00���ŚZ0yr-i��==-e�� <iֱ�T���ir
��R����H�m;͑#1�0jT'V��H۶6�.O���mCh�b֮a�����q��?K�N��.MxA"�uƽ{���%�]�r���R��ti۶={�3{v?�ܚagg&�R"U	�^� 4II����Y�n=Czz.�l�4G1�P�tt4��|=���#F|���gѢAu�K��o�/����r11)�=OXX.�s�Vj8:Zҹ�-�'w�S'[lm�(�\A��d29���l�r���h�41d�Dw|}�amm�����Ό�����og��ws�hk�L�uke�&T�3�ʸ~=��'op��uN��Aff>��zt�l˄	�t�bG���EW1A�:(55��[���ogIIɢO�6���T<=]�UqA)&N�F������||�f��aL���]��#�4����8�ɓ78q�:��٘��ӣ�=��gO{����A�:J.Wp�h[��"((cc=&Lp�׷;-Z�*�<A�ֶ	�v�c��@���]��F���133TviB�0#Ԛ�b)g��$((���h�10Ц[�V̚Տ޽[��d%ƺuFi��	G����|�m;Ö-��s�>={ڳf���&Za�Iaa	w�f���˽{�ܻ�Czz��9��-�,����+.�^*������������ja`����VV&X[�`eU�tC������o����ěon���+6n�J��v�.M� �B��jPjj6!!�Gq�x,��%t�М�����ǁv횋��h۶m����c�e�R�L�<s��pp����7ڶm&Z����{l�x��;/����`,LwZ�4SviuVvv����R�~=��ػܸq��������kӴi#����0��Pmm��ett4��Ѡ�XJaa)���RXXJNN!��瓒�������477��ʄ֭-pt����
GG+���w�Ennl#88��>�ԩ=�]��lsE���B����;GEDD������H����������8w�����.���0c�;XYu%  ���L�6m���+^^���iߠ�l
�ɓ7ذ�!!Q�hф�^��ر]��J�������ܹ��oΜ�YZLMhӦ)���iS��@�f&XX��[=����3IN�"99�[�2�v�.׮�p�vFyNNV�mی�]��ڵe�[�T�P����\y����Y��%��\u�0#T�K�n��e��Lbb&���xz����D�n�D�P�EF&��A``��h��ᄷ�+8ѨQ�����R{�^���D����Z_t݅+H.Wp��m��FXX��Ǔ�W\>���{K:v��ѱ)&&�J�5'��kג��N!**����]KA� �vmI׮v����Y��1+]hh4o����-��i�t,-��]��o"�Uw�������W�};��֞��ۋ��-))���H"8}�
��n����v��ۭ�|�SVV[�����8���1|x^}��Xܲ�22�8z4���h��!##��t��
w��t�lWg&���)���xΟ����8.]�MI�[�&xx8ѿ�=z����#eHHHg�̟HK�a��W�С��K%P9��)��}�}�.������9Çw`ذ��i�T��	����)���h���9|8���"\\���)����L�%
B�$$��a�v�8���:/�܃3z���s�����իw��P�{�V�'�����.�Z��H�x��_���h"#���R�[�V�����urm������ʑ#����)xz�(�$�o"�ϗ�U��]al�~��W�`gg���e-0NNV�.O��R�O���?���H�����6y0��+ݺ�3=	*'""�o�����4on�+��a�w1�9nܸǾ}�ٻ�11w��4���'z�j�����K�q���r�p4�_�ر��
h�ڂ!C�1xp[\]��]b��dr�-���?���O_bʔ�.I(#�dr���'��e�i"���`Ĉ�ߕN�l�]� �y
����D"� **##]��w���Gu�]�Ѐ����o		���Ŋ��=4�����i��w��{/����C��c���t�lנw2��8x�*^%))�-L˃M���D׺�?�'��c޼�,^<�N�\ω0#<*!!��;ϳc�y���pwo���]:�]���$�r�vƃq6�=�D"�g��x{����JӦ��]��@�<y�ի8y��;۱`�'��;)�,���S�޽�ؾ�aa	��2dH[�mO�n�t�y�B��+w8p�*\!!!kk�m�ȑi�N��_��s���1bD��r�hQW.f��?*�_cӦc=���1��ua��.u�o� �uYYG����(((�m�f�����劓���K��BAHH4�|DXX�{;0o�'={�+�4��������8x�* ��eܸ.���uu1�geDE%����D||���Չѣ;Ѣ����{�S�n0s�O���d��i"�(�3Y~~1;v���������������_?Gq%ITDq��'�NPP$��9�haZ����{Kq�$T�\��С�|�M����̼y�t��B٥����Lv�8ώ�u+�N�Z0~�;Çw��Ht�/�b׮���s���|:vl��ѝ>��ʭS�Ą	�i۶~~3�)j�3������	~��,R��1c:3sf1�� �8�\��˷�'������>:���J�~�bP�P!r��ݻ/��7Aܼy�!C�1�'��bR����e�6o>Ahh4��3zt'Əw��5H&�s�h�v]��?��)��;1a�;��;�LKHl�]ƍ[���%�7Ϭ��P�Q"�4$��ű~���"��lĴi����&��:*>>��	����P�O�6xy���劙���KT�B�����|��?7o�cԨN̝;@\�z���|~����r�۷�ӳ�=Ӧ����EeN�������پ�'O^W�@y��=Ǝ]G�����k�1ƵH�������Z��S7pwo�̙}4�MtM�z$##�����:������Z��㊷�[�Y�B����(��ҟ��D�mϢE>�j%^��|�6�7�d��hkk0fL�M�%�C*�aW��;ϓ��N۶6L��ΨQ�����֭Ǝ]��E#�n�%��f곣GcX�:��g���ˁ���[�V�.K�VXX±c�DIFF-[���ㆷ�+;�3��'o��9>//W�yg�X#�1r��������|�6NNVL�֓ѣ;��<U�B����8�n=ÁW��I�M�I��vJ�)11��c�bff���E���!�L}ͪU�����Ñ�����A�d29aa	D��A||��xz����J�>���
����ĉX��i�;��C���.K�H�r��+��&>>��C�1cFo�vm��҄Jx8=�֭��r����L�ދQ�:����;w�3r�w�nm����*�$�<fꓠ�HV�
�ʕ;����K�G���-_��ҥ�hkkҧ��ޮxz���lAB�EF&���
��kז���`�*��T�￟e͚��3=�o�9Pt��.^��O?�`߾���k3iR7^{�o��!�y�#G~G�.vl�8M���,fꃈ�$�-����7��ve�OڶU��AP���\#��ر�R9�:���튏�+vvf�.Q��;w�b���D۶�x������T�ٳq,Y�qqiL��Μ94o��k�U���˶mg���dg��۝7��_kGE%3z�wxz����HĒ5D���,55��??Ȏ��С9˖�k�P%%9r������������)^^.���Ѿ}�J�?U\,%  �A�ڊ�5('��ի��;���	K�c� 7q��������=��yG>�d�X�(.��u�i֮%##���y�����4��c��%0n���߅������(f���b6l8ʺu�����C1�����Z�drΞ�#0�l��[�2��0z0�ƍ^�Z�������Xq���];6n�N�f&�P}�QZ*���8�W�����o�׷��O�k�E��Otu���Ñ�N�%	���T������`���f���̟�Y��S�8���f���{���c5P"��%r��;����)((����3kV?�� 5*::�����ùz5==-<<��re�@g���|20j�w�;���:ZZ|��/���r���B�`ϞK,_����<f�������PL���)˖�f��SL�ދ%K������R[����/!��Y����3{��E���
��7���w��ݩƎ�@�0SWDG'����	Od����� 7�WvY� 40w�fP�bs��u
��-��v��˥|�AVVnn ���H$(
�M����7�B-;¿�:u��>�KDD"��ue�",-��]�J�};�Y�6���ՓD���W�ڵ!����41`���޾Ǝ�fM+Wb��Y��պƎ� �0��JJ��^�ڵ!�kל�+�ѦMSe�%�@nn�_��?���hrr
qv����m>�d?��hh�Ѫ�9~~3h�RL0PQ		�|��"��pd��ab��g�Ŕ)��2fÆ�b2�RR�X�ҟ���ѻ�+V�Tc��%K�`׮0v횇��e��aF��;ǢE;HN�bɒ!L�֫�pAjCi��3gn��A``��DF&�������:j|��8ƌ鬄j���b���?���ٙ�l�1C�s�:u�i�6ѻ���M��B�\��;���͛��;w s���n�2���3"<<����V��!*��+fŊ�l�|�~�Y�bL�̺!�PJJ�8:�GQQ�S��p1c:�|�Kb�c�9F��X��Ń�<�;b��g	���~f��v�Z5Q��!T�T*����r�!����q��%����a�V��/-~q"̨�˗o3{�/����G#y�%q�R��%44�ɓ7��x��P��ڄ�!�M=v�>���1F�2N�������v��O_3|
Uv�n6K��šC�L�҃����A�]pII�bР��ڵ%?�0U�V_�\q�BE(
6l8ʈ�Ҫ�G��+�� uR@@���x�J�$&f2`�J���pW��RSsx�_>����|���ǈ S��)��ʏL�ԍ��ǈ�C�4mڈM���n����w��Wr��jۿ��1~~3�`��j�oC%ZfT@ff>�Nhh�3��_�/��P�,]��O?� K��=�@�P �(P(@"��O	e��>�))I���U��AW��\��9FQQ��8U��g�ҵkWe��D))Y�nn���2]˴��)))Qv*�����O>QvO���˻����?�i�z��êm,�o����w��O3��r��}6@sŨ8%K`��_ �믹t�l��A*/>>MMM�n��G���������hjJ���,��    IDATPCGG�D������� 45%hi����N�V=���(�T*G� MMe��q��q���3��2f��K�F|���*d JJJ9r$�&MRv)*��ח��xe��Lff����`��,Y�'�O�`ݺ�qt|���&N�Fdd2��me���88��j�B�%Z��˗���Éի'bb"���|kք`cӘ���Vj!��cǖ	BmX�|?))Y-RɁ����l�w�Vv	6rdG�t��7�0x�*���L�������� &&�i����##�j��aQ�KHi����g;�~������?�AF�PTT�����3�ڵ��+p�v����	�bӦc|��d���]�� X[���o���Y��/f������ڧ��:��O��TƼy���6��|"�Բ��|&L��.�e�k̚�O��Ae�����U����{�O�8q=AA�O\7Fj[zzl����ӻ����uu5������^M���k""�^h����_?�Ç�Y��H�ڀ�nf��ƍ{L��@�"�+��-|�vNNQ�G"�F�t�O�R�
���-�ʀ�io����̀��{1qb7,,��Q� �t���5aѢA�.Eh���[�^�W�[�g��e����+��ɖ>�G�S�t�ڲ���D��%G��0k��89Y��7CL�)���_B~~1���� ����+F*���_�T*'7����_�LA^^2����"
99�BH!
�-k�W( ;�������Q#���ut4���x�~mm��u���}���.��F�t��P��@M��504�ASSCCm��5�����@MMu

3=l�IK����� ��]�6�={���/A� 00�C��	|[,"*(���>[���W_��[�s��->�xZZU;��9�7g��1{�/����A5W\?�0S~��,��ॗ:���*5�VTUq����|23��*���/&?����Brr��.������

�˃KNNQy y��'��ƺ�I�ɺ������Ʀ1jjuQW�`h�S�--�G���{jͲ������ꖗW���9?���R�#����WR"���l�ל�"�r��R

��+z
��IM�)ߧT*''��TFnn1�ť�����&00���bee���!�Z�Uj?�����v�-�����k�)T���"�}����Mѻ�I��u�2���|�u��j,^<����[��L��oF�Z�%	_}5��x�-l���J�Ч�D��a6壏��x�`����r�_JKeI>YY����}��df�=v�~~ypyx"�O��Z��k���M�Fz��ka`����-Z�bd���^��e��-���@��tPS�<�2!T���^�م�A�a�����Y�&�B��J�H$��� ]�ͫ�kޓ�3\ԕ�QSu֕����Z@�F���y��^{�g�M�Y>��*�u}�k�I����V���Kxz����Ӧ�1x�*6o~WW�J���H���1t�j֮� �L��KV�d��1L��p�Nj_i����<RSsHK�%##���,���HO�%55���<RS��5F��Pcc=7���Xcc=Z��(���D�����VSS�x��������Sff> �~����T*GCCw�������FtueO�F^ԍ���;ζm�k��CBB: [����ObnnĘ1�=���V�V���lm��w�|^�F���o��Đ!�*�k>�`8~��^�Zӱc����a�(
>�`��z�5k&3rdGe�$����$&fr�n6ii���咚�MFF���RR22��cd����M�`nn��[3�͍033|$�<%�zÕ�_������0#����:��2LM��v��Ӆ^�Z��_�BB�W��O����ᇷ>��W�����Ӷ��������cOz�I����ǯx?��'ݮ�~�U_e�f�ҿ2��R�hiiiPR"�޽6n<ʺu��ٙ1vlgF�숭m�>��ݻ����q����ό�tؼ�>�x/����E�|�?߳ҭyӧ��ȑk̝������/B	�&�L5��������w�M�����쒄:B*�s�^II�$&f���Irr��og����|���ZXX�SSZ�6�[����ann���!���055@[[�Յ�)�&G]]������7<=]pq���.6�����	ӳ�������*z����U����~���?����_��R �ǳ�ǧ�jU _|q7�f�ۅa��Wy�De_w�zm=�"����j���X�l$MY������/�Vj����3�d��?Y�zRV\��3�j$�ʙ3���a˖���C��#�-'��<�$&f���ERR&IIY$&��޽�Ҳ����XY�`mm���1m�6���++c��L��lT~E\���y�IؠAn�N5:�Nm��T�X��Z]�ǫ���"���l��nȕ+�14�\�㾈�R9˖���˕���k��ec�a���H$::�e�v��j��A�*�E^w�\M�d�mҤn4mڈ�^����<֯�R��e��Y�j"/��'F��P���]�x�U�L�o�ʑ#1l�>�v�l�]������NBB����ǧ���N\\�#�*FXYcmm���166��o[Y�լ�:�����[�Vx���r<���Ue ����c<�����T�Ū���,zzN�Tz����Ś��S˻�=�DR6<��w`��)ܮj��������럪�w�.�x�/���֭-ؼyf�'���w�c�yBBammRCU�YsE�L5���,\�G�\���E���X��Ӊ�K+_�D__[�&��5�g��L�ܝ�͛`mm���q����j��ܳ�Q��^cӦ�4����ܽ�MϞ�Y�v2>>n�~|�5kB��K��<K���2��Νm;�S��GWׯ��P�ג*�Pu�؂={�1i�zF�Zöm�hڴQ����a?�����~��R��qF��
o���p�m�E��͕]�P

J����͛���O���{$$�����ҫWk^~�;��f��5��)AjFm�	eLc[_BRE|��^�v�SZ�yu�RNN��ۅ#�cii��/W}��睬��k@j�K���ٻw>�&����߰m�l���+�����VMd��o����b��ǈ0�
Ｓ��{/�u�kt�l�쒄J*-�q�z*11w�v-�����Ĥp��}
�#��wo�L遭��Z�cn.��	zZ����x|���c?��;��N��z���[]�Up�l��_!0�me��MͲ��ll3n\F��H�V;)}���=���2���u�T���!kڴ�v�e�T?F���_}���.�oߜ�s���{�۷-Z��p�u�3/��v��al��
ݺ�Rv9�3�drn�� ::�A`)/��iH�r��5h��GGK&O���4Vv�PoUu���'e���Ek��c��:�[��*�L����)SzҦMSe�S>^��Ԁ1cʦb��.�5�ڪ��j��Ր5j����f��_7n6L��
m�p������o����X��f�h͚~���7�B�^��]��w��'66�kג�C���K��P���GGKF��@�6Mqr��E�JM�(� Ԝ͛O���ŢEʟx`� gn�Heܸ�t�֪�N E���CGG?��,^��������)����ij����5?�x�W^�Sժ>f�`��|����֗~��]N�%�ɉ�K#""���;DD$q�j"99�H$�7o��CS<<��3�?m�4�uk�Z]9Z���5�dR����X�� ˗���������ɲV��ݸuu5��r::̙�K������{��g��q�Y31��3��ҥ����=����i0�R911)��'�Dxx�|����hkk��h��[3�k���5m�4���D�$Q�-Y�:�`̘���RW��f�"�H���(
������2h��'�x�́��s�����_~y�*Um"�T�ŋ��3�W���`�e�S�ݾ���˷�t��+<<������qq��m�f��v�ͭ�hmA�'��+���c	],���D§����ٛ+h45���q������0th��(Ue�0SA		�L���A��X�d��˩W��
�x��.��ʕ�𒑑���:��Vt�МI��Ѿ���b�� B=����{��ɢE���m��r HM�毿.bh����6zzZ��iad����߷+�� �SU��{K&Lp�vѷouj�T�$�Ldd�1i�89Y�j�Dq���ťq�B.�s�B��wQ(�ֶ	:4g�Oڷo���5���%*�P��dr��ߊ��5�f�Sv9�#��㽨���Pȑ˟�\mmtt4���"%%��W�P�U%�,]:���>��@���8S|��R3f�����6�ݙ*��D�իw�p����q�|<y��hҮ���.���P:w���X\�������\����&T���&**���E*��޻�P����XJq������Hk�2�>�l�11�gٲ̟��1c�СC�\�]���X�x7o�c��5�&��*)�r��-N�����7�p!���R��qwoży���7�f"
B=�m�6
��9cU~�D�@M����)PW�#��������) 	R)�i����ݐ>|��??�ڵ���2Vv9���mB�Vfܼ�V��kj�����w����邯�v���������4�J�iܸ�ϫ�v��ɤI5?S\]�x�ٴi:��.O}��ѝؾ�<���С���hx�L�0���᯿�غu����U5��ɓ78{�fyx��iL��X�bݺ�+�
B=7a�JKK��ٓ ��L��j��.b�� �4uuYM�*T҄	�߿��;..�9s63sfo��P#�xQ����PZ��ץ���n�Z��w�177dɒ%ܸq��q�TBA�yy���i���Ea�ߧa�z%��Ϡ�Ǝ˄	�]��yh�R9�g��/��JϞ�O}�矏��/ظ�h���J�� >Qppӧ���/1eJe��2d29��?��㱜?Oq�����aO���t��
���.U%y睝������=��&�C�l�0KKպ2/Ԝ��"����M���WUn��[�2	��?�s��>��J����ʬY}�H$��r���^M$<<������P(hj�#�+t]� 
��_@ǎ-j�G��LάY�9q"�]����d���ZȺu�>�NC[{f�3Op�Z
#G~�K/un��JHH//'N\'+� �F���@�^����k����BC��<y#���<NMM�B���,\�� �G4T��%���FRR�9t�-���-��9>���(��"�~=##z�v 4���%��F]]�f�Lذa������Ϝ={�|܌��r���cn$	�}�+֭���T���DG��o����*)����%��Mؼ��Z�R�D�y\NN�}���	��6K�Ն��"��������֭�����Þ޽��ہ6m�*�LAT�\����x&N\OQQ�S�������6��O�W�ֵX��l��2�N�DTT�w�Sj7BC�	
��ȑ����3��ә�]pwo���:s��W�J�B�D"A�P0~�;�~:==-
Kh��
[MM����?�5��	�DNN�&����|v횋�E�'>��雌�?����<��zB��R(���O\��H@�h�X_�%՚k�R�&44�s��P(�}����ۆ޽�ر��/�K9q�:�E���C�-�z���H��I��Þu�Ф��*���T�+���ŋ�ع�u��m��DG�Eppaa	��Ipwo���.xz:cgg��mv�țonA.W������&�WO`ȐG+ܼ�$��'r��O�44�:�=k�N�=���ǰaߠ��ɮ]�ښ9w�.^�ő#� �Ƌ0�O�օ���ٽ{^��ޮ���'����׸s�>��xx82p�3}��S%��TYYG����(((�m�f������JTT��m�1e-�
�}w���_��50%%R���±c������X��q����<y���HBB��?�tf���ϻ�us��*���} �t�cݺ��ؽZ&�3`�Jn޼�Ԯe길X�w�|q�P����,�������,tu������L����E�1{v��/���0�Й37;v<�i�z*�����C``���:u�����<0.�kg�R����Zn�� 00���pΞ�C"�гgk��]��v�iӿ�>de���A�	���:���l�4�N��@�&+��3~$::��[_����))Y��D������b���.�L���+�y��;177b�|�gvA?z4�I�~�I�W���4mj���[���VI��S;v-�;���7���ŕ+��w��'�k�3f��$���Kz�r`͚��.�Zݸq���p��ùt�6::���爧�N��*�DAT�B� <<���"��J��H������q���Cç_�1�[Ο�G"����·�N��H�Aܺ����(-��믯Һ�E�C.Wp��m����$22Mz�vx��T+3�>|�%K��������Gf�SS����ɁŸS�\�x��c�1n\V�������k��.|��X%TX�D��J�����\��&�����C��	�ƍ{����劏�+�{;�����2APQ��2N����8���$'gammR�7�[�V���O'x��?����L�޻�+TQX�-�O߄�Mc~���̪�ZNNǎŔ�����Ʀ181p�={�F[�v����l�n��+�a��3w� F����I0��%���1�P-#�9�'�{o�זپ��m'0�m��M�E"̬Xq�<���[�je��r�D�Pp�B��]f��+ܽ�M��䆷��;�6�Y�A����BBC�����ȑhrr�pq����//W�ܚUi�r����R����E"��
?�p�+�3`�3k�L���A||AAe�/g��!�+��ɶ|�˳��	
��;���G{���dŊ1嫵�Y��D&�#�HX��%�N�����x��󛎗��#���
�Y�����6[I֊�fN���ĉ������U��T�B��ҥ���w�}�.���E��ޞ�����tAꖤ��c�"8s�&
��n����v��ۭ�-�&T���\����ɓ�Y�xs����x��Rg��IPP��i�ѷo<=]���Ii��$$��x�NN�����y��h�?^R"��e)���̞ݏ��w�R��%K�`ǎ�����o���Ug��1j�w���k�T~NNׯ�֗�7�ܿ�π+�޽�ֽ��r*�ʕ;��Ν��liưa�>��0� <Sdd��F�������_53
/�ȑk̟�}}m֮}�J3�fd�EHHǎŐ�S��CStf�@g:w�S��R���eժ@���X�r�S'4�t�6��Q,X�%zH5�ᢚ7o����GƆEG�������=����R~��˗� 6��Gx�0ÌB�`�4?bc���3�����Lv�8�Ν�IHH�ֶ	C��cĈ�6�� u�T*�̙��@���IӦ��g�ٳ��V����,_~�m��0jTGV�S��V�BAdd2���Gq��m45��֭^^.�L��5�T�իwX��w���X�Ћٳ=�{HP���"F���ݻ�ah�î]Y�`��2�����r�ԩ�����2�gg+e�^f�����|���^O��Dʾ}�ٱ�<'O^�qc}F���ȑ�Ռ(��P^^1�GAHH4��89Y>��F۶���.B�y8f������·�d���ݮ�����c��D�����������퀾��\1���Y��_е�_|1k
��ܺ��С��ر66����1$	
��A7O	r��kI$�aô-�Z�mK��STT2}��ŋ�d�IJ�d��l�v���"��w��o��;��?� <Qjj6������s��d29��-Y��ooWZ�P���B��%p�bS��bѢA�\|�Ν��~������k���vc�@g��T3h'$�3o�6�����{Cy�վbM6A�haʪUY�l7��� �k��
�ѶMMu�k��Ѡ�Li��7��B�.�̙�_��<���8~��AA���2cFo&O�!ց�bb�>X�%�˗[9S�    IDAT���ʕ�8�}e�(�S99��Z���1ڶ�����pu�w�g�LNXXB���������۷˗�Ā.*��m��-�M��:�V}��V��Ν�c��mdg�ݍ�Y�r�ne�Be5�A���+q��}~�����"�+
�d��P.\��ݽ%k׾̠An�F�G�drΟ�/��,!!33C��\Y���>}��ښB�TTT6xx͚$��ӗ������iVVG��Ihh4YY��6a� g�����a_'>����X�h;AA�̞���Ń���/A5��cٲ=(��0�'�ʹ~�nWV;�;3,,��?�ʕ㰱i��Zd29��ڵ�ܸ����{�Σsg;��%�j),,�ȑ#
����|���2�>>�t��B%.���T*�?����de��+}x����p�z*AA���Dq�|< ]��d��xy�bo_��p
��������A�n��]� <աC�|���*mW?��5�	 

J���{{s6o~Eiu��
����_p�V:/�ԙ9s<pph���AP-��y���?KI��N�l��.�߲�t,��B���~���{L�ԍ��11������֭7����	OOg��s,:uIaa	���n�l9�ر]���*?۩ ����;ٽ�ɣ���G"�����N��>CØ�����d��K>��R��*
���W_p��=F���[oyckۤ�kA��ť��N@@aa	hiiл�>>�xz�Ҥ���K�Lξ}�Y���;�����w�[J't/蠋B�,�e}A�d;@���DAd�Y2E���@�m)��N(�t�M~��N�H��y���朓�}Ҿ�9��凉�Hd��L�֝k��~�"''���%8ؗ�@W��r�f
Ӧm 99��>��A_�I�e�<y�7�����
�.h�OO�:���i�b���(F�Z�ʕ<�m���\���&,,�!C	퇻�f���j��䄅�����7R��jBp�}��ӣG+���m�@�(((d۶3|��Q���ӵ���V\�ǥKw04ԣK������GGKu������9���e����hyyR���wV�:
�PTT���l�8��`��7��h�b������GV��X�s�ǧ�h�~��	�sgw��Za��@���r��5����W�{77�f���O߾��o�B��l4���|6m:���Ǹ_�����Mjj���һ�/]�z6*�-��p�>֬9ΤI����!"�_�(�r%�Y���X� ���r�\Y�Y__�>�ԩϨ�TUи��|�����p���6gNN>˗fժc�ٙ�v�$h]o���CZZ����W8v,��\)m�:3e�3���O�V"_N�>n�H�����Jwpe29�����{����8o¥�?`ʔ�t�+V�g�� u�$�G~�=�5k���g�!�ˑJ���d铟_�4�ok~�F+fΟ�a��|��zɓ������>��7rs����@�L��IU����Ĥ��W8x�
��{]]�t�����o_?lm��m�@�)((b��#���?ܹ��12ң_??��kM�^>X[7��7R�0a2���{_��G�4>��tx��@h�O����r	yyR����H�Eܺ��nSkM�3�J���o1��f���Ku>߹sѼ��"#		�̜9��ROú����;w�enM��ɉΝ;�ی:#..���G�fh��ĩSI$&>��X??K��-��ǟ^���ۼ�X��Czz>�6����Ld29&&���̈́	]x�i���#��ĉk���&<=m���ɢ����PXX�޽{���R]�r9��w��;o��W����Φ9� ��_?��9�J��g�����r�Q�y�N{�de��駿�q�)�v�⣏���̲D"zNT�F���L�<���׫���I�@tu��ϿI~~<�Lc^g�E���A"���z8���X�h]�z�ۤzgǎ����Đ!�,^<J�����Æ��9ttLh�l���dd�¢/Τ����yUI��Ɨ3s�f
˖b���u*d~��2ｷ����K�2|�Su6WuٲecǎU���[�2n�8u�Q����3v�X�l٢nS�mXg�E���C"���[�RȬ\y����k}x��Ɵ�����@]7�֪a����i�3ﾻ�V��4�k������{����߯0|�S̛�,���	)�@P9r��E���r�Q,���"�S hl4*1�k�9N������T^�T&��i�i>�t?VV����Kt�}w��@ ��r9ｷ��[���o��쳁�6I ��F�df�2�&Lx��m]T:���w�5�G��bx饞��F?���U:�@ � ��y���l�v�u�&ӧ���MuD�3�~�+	����T6�\.g����=xx������8�l|�@ �E.���?�s�Y֯�B�^>�6I �!�B�\�ǦM���q���d���LBC�ĉk̜هٳ�j}��D��Ĵ�Y��)*C5�b=��j��r�?�o���a׮s�_?�=��m�@���{���ʊf4��W�/,/�����_h߾Æ���������snݺ��ݯ��[�^�@�lu��TgL�\� >4���o����n3JQ�A��df�r�|2Y�Fˮ��kQSכ����X��0�ןd��	B��P���밒?�K�=3{�^��������Z�A33�;w';w�#$�3~�,&&*�T ��/�aذe ܖ�oGϞ>B`k֜`��߱�6e��6,�� gu�%�"6n<�'���ҥc���_���zB��Lnn�cԨ��>i�>}�Y��RPP�ƍS�&Y���QQW�}%����U��%�kc����(?p���_�IC���ѹ�;::��3�P���������}^Ѿ��VE�[���|)	��f�n�_�Zugg+F�l�СA��ۨd�ʾJ���vVLu���Y����}��-�b�ٷ�s�����1bD{u�#�%�eU���y������*�j�F���+������o��2������%K��_?>�|$VV��7������U�u�=�Ve�����(,Tt����gǎ�����w}6P%��Խ7u^T�}T��j�Z�	��z��RXX@\�}��������#F���g�booQ�9�����j���κ�ɾ�.B�Z�'O^g��x�垼�J/u�#���i���ME���=�WW�a+f�Y��0�����iZ�1�����W��o��GC�4I;�i=n1�t_]�"(�T��`LM����w��5Jq'���{=�t����[���>��&""��?�ς{i�ލ���3hP5[W3���jr\}���\�|���2rd�}Wu�LM���+��`��ye���|5Ec�����5c��gj��S�n0c�&��س�5ڴ��چ��?/��Q�f<�����xL���s�>�|�'���СCj[��Pu2�����r�z���+���Es��m�z�g�ѩӽ�7�!�����9B�lc!11���ѵ��~:\�m�\Nbb5�@�
U&��Y�lβbK��̹s1��K��M���zo�dX���|��H��s:_���w�������ou��5#33�����ۛ��w���_v����C���Z�͍��ѝN��y�)W��}�Z[�����p��FEhu��\.���o]�xп�j�655��3EXYY�5����+�Z����x"g���ԩe�=F__���T������ͧ��"T�ДuV[>�x?k����t(*��
3�1cZ��X΢�k��Uv��f�x�卤��u�K�����C�`����С�=�TZ���.���t��I��n�k熵����}�w�:��5́�.'f�o?˥Kw���9�z]XX,S�|����++CEU�jK].ںtUj�F� �z�m<pY{J�[�ں�T���.��E��ث� @1�I�/������qǖ�l=.aW��ʙ;w��E�{�k�ښ���������e292�"�����b	O`Ŋ�����dI�.�t�ؒ���j����'}���\��-f����>��WBB:��m_����ӿ����v���oC077�C+5��N��=�ξ��[�����;�uU�������&�{�=U�CP���B�������P��
U'�V�Rپ'�K�˳|�a�l���[_�ǧ��A}��`��������Ic�γl�v 3�՞�&�njrn��XO�W4J̬[���y������Ri���ٴ�4��ڛ����>���)B1`@�h�)h��#�#�f
�]����'�����ӵ�������w���t�066(�#��(�Kmm��|9�Z�p#f23s���#L�ރf͞c���Ŵi�	O`�����4�hnnӦ����OO[���pv����J�\���Ѻ��6M�sgw�41T�9�B���˴i�бc�~�S�n�u��9y�:�g�Ȍ�x�.�6G�E��rRR2�s'���t���HHH(^����(�755����bF__�LΰaA̚���ɸqնM��j���H$��=�x���1L��cc��E�Vvuo�
�͕r�H$�H$+,,B&S,P}}]-qs��ͭNNVJ���lU��z�k�K����[/�� �)ff�t��n3j�X����D�N����ۋ^2�S�UIHx$T��I��Ŷ��te�]]�7o���t��
GGK��?���0z�w$'gV8���.	��43f���Q����5�_|i���{7�5k����h������y���mt��ɷߎ�Ȳ�VVMpp� !!�Tl%(B碣�}}�H$��"�b���E~�Lf�@�R�		YM�N|��QNP-yU	������E����G^�&Mqr����[�w����B)^��̫���d��,FOO}}]&M�Ƌ/��y�5|�G#��ҥbff��ɕ�R���|���,]�'/�ܓ���q�%�С��]���raR|� �M��Fbhؾ>L���HK��d�E&����All*qq����Ollj)�R|���#���''+-x�V8:Z<|n�����
D98X �+����t022��{0eJ7,,D*U���Lll*?�p�E����H��c��̞�#��v�/��ر���J�Ӷ�+��_|�q:: �K��Ń�?I�́�uo�@ uDffcƬ"7W��?�"z�h1w�fw��X)/Z�Ŋ����V��X��nC�n^�0GG�*{UT���EEr,-M�9���?���f�6d������qr�b���OI�bҤ�ܺu�-[�kl�v||���CXX,.�QX��p1]]],-M����4Hs
�@PYYy������ٽ�U�64<23s����,11�ܹ�+������zz:��[<,�t��gg+\]�qq���Ƭ��!��m02ҧo_����Ӡ�����u�+ƣ�W޽}�#V``�ǯ�΢e��j���df�q�R,���RR������ˎ�@�{�ｷ��03==]�rӦu#4���W�� Bf5$$d�s�er�@s�˓*�I\\i�J\\���ښ��(hԿk\]����-+�l���0xp[u��5H�e� �9s��+���7��f�����u����M�v%;�d��*�����p�BU��X��""#Ky]n�LA&���`A`�+��.�����#Wzp�\�_b4	��� 7>�|d���]	M�1W�<y2�ׯW�j��؇��[�d��6�Q��ڢ�봾�H���ĸq�x�Ѹ�5S�I�HO��1+II�b��W4���#�)��=+%�����Rki�D�M)n9Q����U��bܻ�ͬY[�7�33sKs���/U ++�LFb��,sb��:��Ĥ��^��n��9�
Χ3˭�7n ��փIU%�	��Wi�E�q���ڛ�bcS	�%,,���c�r�yyR�65�Mg��oMP�+mۺ<�gL�-��JB*-B__#��ʈOU*ZN�>͝;w��5:����mB�2�|�n3�Bnn!�~z]^~�3�����ƾ�j�6���$==�={b9x0�;��nCp�/�z�ҩ����x߽����ߑ�S���3qq�V�=��de��������11�DG�%11CEҤ�!..
�Ҷ��>�*..�Z�7r�B,G�D�赁�����Ulܽ�Ƕm7�~]!�~�i�Fɪ�|Z��ѣG]٢6N�<���22<.�\����1��f������=AA��׉�@<<l��p]Y�^a��ѝx��=��F�Νk�~�ggg����{�^�=�;֭�Ͷm/ר�����uZ�L���2Μ�ő#<x��+�affD�����K�^>���r�f
�ǯAOO�_~y;;�z�_��޽l����Jt�#��ʽ{ـ�"���nnָ�6�g�JyVD~t��
c��s�t���::��j�=�N����I���?Y����O�ޝQ���tu����zB*-�ʕx.\�Q
�[��"��qv�"0Е�3{�B@�s��תC�^><�\;�N}��m]T�.���ɒݻ_%$d5C�|͏?���w��L�@������=x�i��Lt�=�Сp���FQ���@W������??�:���o2e��xxزa������|ڌ\.'!!�۷��<z��Q�������b���5mڸ��A��5�ͭ..V�K�ǡ����Ϸg��S���*BOOss6n�JP��J�8x�
Ｓ�{��J�_����w�˙ٺu+�ƍ��ѣ격�X�p!���lٲ��FG�{��Hп|9���B�̌�(r]ڶu���LVV'�%""�͛�Ӯ�jOAc!''��ǯq�p�_%%%{{��}��ۗ�]=UZ"y���x�͟��ϟo��(�%))Yܾ}�[�R�}��n�}��B~�"w�iS#\\�iѢ��͔�7�f88XhdRC�ʕx����������m����Tꍌ�M��vr�h$��(r���m8q����@(�3�����p�|l)�KZZ�����:�ʄ	]t�ݽ�H�4��M�ز�E^zi�F�`��I���n��G�&������r.^�Szm6o�CC=�t� 8؟޽}j\iL*-b��=�_�3z�����j����H��͛w���DG�#+KQ��؀-�Ѳesz��a�����Ь����3ٳ'�m����̘���
���H���X�t�J"y@�Z��0K����S���0fL�(�j��3cccGh袇���%:� nn�h�VQY,0�'q�H h$���_~9ϲe!"�f
U%%%�C��r�p8'ND������}���K`�+��O."������	O`����s�


�y3�7R�y3E)^nݺGZZ�iru��eK�ݛ��+-Z(<,��'/O���Wؾ�?��F�&���.�7�]*ԬX����@^}���D����x�͟ILL���(Թs�X|J�\�LϞ=k$�._6c��XX�(�����X]��񢧧�ҥc��0aƌͤ�f1iR7u�%h66M;�c�v"?�������Wٳ'�e�aeՄ�=}��Go�̌ˍq��5^}M��믳��S�;ixܽ�����ܺu��7S��J�֭����G&�������-Z4�M�{�)����ѲJ"R�Z�r9g��f�γ��FNN=z�bŊ��ad�Orr&7�R�FWW}}]V�O���UbG~~!�?�-��G���S����աK��(d -, вe6{�ΧEQ�^ �6$	���y�̝�����"TCC=�woE��X��9���8tH�6s� t�В޽}	���ي�?��ڵ'2�-�>��M���.������T�_O��M��E��]e�HSSC��m��C�����<�i.�����ص�;v�%:�>>���F�*�?mkkF׮����u��th�̔~�������IJ����h�J�(���э3��P̘�	!#h93g���֌9s����ɗ_�B__W�f	���^^v��J/��p��5���*˖b����^y�'o�5�Q�rr�~=�kג�~=�7R�q#���T
eH$-pw��m[F�h�P�؈�����<����g���[4kfʰaA�ձ���%=�#'NDѺ�7NUy�jWWk��#������bC    IDAT��=��z���>����tJ�Lq�W�Я�={*��+V�5��}]�1c>�@ �_F�h���S�����,֬����,j���	�>���|���|�͟X[�Ҥ�!�~{�N=�i�C�^���hf5в��ڵD����s'�\���>6�liðaAxx�*�,��'���d;v�]��r��e ���شi=z��rh���m14ԧO�:�[;��o��k�z����=4���بם�<3�����t�ʄ�@ Ԕ��[�s�Ə_���߲i�4Qj] �%�����ۈ�I���3u�3���w�Ç#8t�*ﾻ���� g���O_Z�vjp!��DTT���$�]KR�CC=<=m���%$�3���x{���l%rY4���D�o?���a��d��Sn|��0�	�̬�����:�����acӔy�e����I-UAM*-b����[�$*3��Te����@ �����:cƬT6�tsk�n��#''�O>��Nҵ���O���Z���ي��0qbrs��(
g˖���߱�5�wo����ͫ^=��\��č)\�_N����%DKc�޽lv�:�Νg�|���֌ۑ#�k̹ ""���ѱcKƍ��'��=f����ԩ��-�[�.gF ���j;}�3a���͛�Ѷ����4�L��?���~#?��ŋG3rd��zY����ן�}����\����CW9t(��~�}}]:ur�o_?z����źұ�Krr�ቄ��s�j���ܸ�����w��C!Z<<l�����QPP�\aǎ�;���>�a���t�ز�yGbb:!!�qwo�wߍ��� oo{^|q0ztG�z?5A��Lx�&��iS��?�XXӴ�1ffF%�kQ h�֦l�>�_����߲j�Dz��Q�YA����̛������tfΜ�ns �H��w��ߑY�����͡C�>�g���������N���S-��{���J��v-���""�zU񘚚���������ˬY���8ТE�*�-�LΝ�f۶3�����<�wo�W_�a�� �5��O23�	Y���1�6MS�����Áo0w�.n����N�aeՄ��<���"33���df摕�[.q�ss��133V�����1�4mjXJ ����b���cbb���Sy��mL����c��.�6K hpDG�c���8p��=�Y�<De}c��M5��Fu@*-��oq��U�̊G��0�{�V�ѫ�&ܿ�Õ+w�r%������y3��CC=�����u 8�����0Q����M||?��;v�������3sfo�����[AN*-b���IO�e�����D���e۶��d]�R'b�lNK�<��滨*O�E��.[��
���#++���\�cFF��y��II����de�"��ˍ��#)�*��)�233��ܸ���cLLo%
�������W_��E����N�����CD��@ ��d�|�!6n<E��ٲ�Ez�������u��Փ�]=�7o(�o��_������L���� �ٙ��cO�޾��Z||pw��-#''���/�m�Μ���U�k��Ϸ# �Y����\���?r�R�w������MR+*3%�?.���}e�?�y]`bb���A������C
�O���###�;w�J���[�E1zz:%NY!�x455R�W����5э*���^냫�5�fm%.�>˖��
����,���0�6����>Ƹq��\$$'gr��.]��ҥ;\�|���t ,��5G*-$6�>��������jM���t�≡���h-EE2N����mg��K�dr������'ӳ�O��o��'��o��ly�n����?x�GrrF���41�I�Z5�*�R���������!::��kr���"��u��G?��ϙ��NM����@kx��@,�4iÇˆS5�/�@P���fŊ�l�x33c�!!O��y ))��h�t)���L@Q��uk'&M�J��N8ai�(�F&�ˡCW9|8�Nall@�n^�һ�o���۶���HƘ1�?�ZS��Jb�����q���ڵsc޼�ҶQ�~��Q���˖��kWOu�� ��˸ �n�ʸq�ecʅ��؊�4,h�΍�@W��\pnt^����R^���8t�����+��@������d�P�8z�I2V���t�D�����GH�j��ټy���N��q�������ٸ����̜ه���*;Ofd< ,,�b	����XRR��H$��Z�D@�3N�n턹y�.J�9t(�C��9y�:yyR����O?ڴqFG�����a6 �<�Ųe!�U!55��{�ض�?.]���ђ�#���s�pw�Q�yu��ͧy�,X0�ɓ��ۜ��L�3��v̜��?��IM�F__��\
r#(ȕ-�i���\^�TR���b1Tڃ�H���W8���~��8�rEʆϕ,� b��Iz��L���W�Y�j"ݻ�R�I�ʉ�H`ժc��}KK^y�7&<]+��'���x��b	��8n߾���%mۺж�mڸк���+���r��u���Ν4�53U��y�V4mZ~���{<��"@�`jjȲe!��%�����B����p�HzԆ#�ө�{�ĩ&�{�y^{ms����׃�mNCB�Č��-[�l)�=&&���Ν�!,,�+W�)((��� W��\�����v��ddgG(]T��1;;�\����(7��±MLʕ�.���
�Ǖ�+.��ؿ��E*-�7~bϞ�|��Ǝ�n��Z#��9~��}w������Ǟ��{0lX�'+*���ŋ
����1\���TZ���	��.J�Ҷ��Z<�ʞ6��Ǡ�#�cGw���o_?e��u�N0�e�S	r9L�܍>\��f�;î]�ؽ����t��ɨQ�߿���1<x�i�60mZw���nsB�TDAA!�/�s�|4aa�/���T$	���	
r�m[W�z�oo{�!�c
e�
(�����RT�{Pn^��±MMˈ��KU()���hr��%K�d���rO�{o���$7��_~9�ڵ'��H�[7/^~�'ݻ��rTBRR��Es�|aa�\�|���|���i��I)Z]d7���������?~����lٜ�`?����.ŕ�P���C˖�Y�f���j��q�Ʈ]�ؾ�?n�H��ÆQ�:���O�*Y9y�:!!�=��|2\�#�*A���r�naa�/�s碹p!���|��pRzpڴq��ɲ������R��^���E���ۋK���קl�\q���+�4��;����=�Y�,D��hׯ'�i�i�o?C^^!C�2}z|}����B._���YE�ٳ�$&�������-mۺ�.�Ziލ��B��w�Ç����+DG߭�����.::.|�����li�$''�_��Νg9u�:��&ĨQ�E9�p�|#F�`���|��8q�b���)2����$ex���1\��LQ�kkSڴq& ��6m?�v'�1��_X.N!xr�y����r��Ң
�.[j�de��M�JT�{$��G�	ꟳgo3e�z��MY�~
����6I ����.�i�iN�����5��?ͨQ��6��5����?�-.(�.Ri�֦�x�ڹѶ�K����]ॗ6U�&�$	��ך%KF7��Yu�L&�ԩ���y�_��TZDϞތݑ^�W9�����a���Ƀu�&�^g�S���ѣ��l�;�;�رcU"f*"''�a9�;\��ŋqܾ}�\������,�����}����,���[��\��s%=EEE�r�J$�RWK������Kz��4i\#�Ebb:'�#>>�U�&ҥ���Mjp$%%1{�l��*�����dg`e���]6���Vqs�`���%�K))Y������H�vn�Ю�[�S5����_~9_������bii�w�M 55�͛7׃����W�IK3�i����X������m��	O`Ԩ���q`˖�Z-�@y1�PO:��beUq��2~�x�����<._V��K��x1���T@�𫤸i�ƹT�|��"rr���.n�ZZ�<���=J�©�����:��@���*/�]���X;�1˒�[���?r��e>�h/��E�&5(�o��1Bݦh-�b`P�ܾ}�v�4	�̬;vv����S-�N7��OB&����>���k���rh֬�˗W��^E2200�cl,e���lٲ��cǪ�,�r�J<�G���#6L���j5(/f*�fm�رH�}[�/���p�b�R�\�G|| ��V��M@��ȩ������#AT���ƭ�dd<�p�⦬
QdR�+T�X\PAQUΤ�~Mm�*����C|��Ə�̂ω�i)3r��:�n����S�����Q�|^�G��K�H$�ϰ\.G&�W�/K�wٺ���6��!�H�^�\����+i�օu�&	!S5fj�U���C����}w'+WNP�9�����[��Sq�^v)q�v�_$'g(�)č��֎B�j���!����ע�ci��x,�ee�>,ǭ�~�^�n�-�?3�b/���n)qS��v�
e�I�(�*�Hx��`Z����W�p�F
�WO��J�o���,W��������@��`nn���!&&��`aa�����33#LL14�cܸq�6_�����2f�J�zʍu�&k�=u�1)ss/Ÿq�4���Q�I*�Y3Sz��)Ռ+99����e��#��d��b���~~���;���(ND�zEnf��c�Ǩ��vI�S|Lrr7n��P��7e54�+W��j�\M�*���f��י4i���W|��||j��ə�9s�~��E�A��IC~S�f��s�7n;��v�$�կ&u&��Û�c;��;��رe�O���5#8؏�`?嶤��\���U�ώgY���r9&��;��9~~�xx�j\yL��`nnR�^=2����lϡ��s		�%r��<xPqSVcc�R�SӒU�*�333��ޜ}�^祗62d��,_B�~�5~��N���bff���]�0�i����m�@ h$g��b��5t��ɪU/!S4J� |�᳜8q�w��κu��mN�cgg���9}��*�ee���ի�\�ϩS7X��/��"���������Q�J�(�ё�Z����+SU�����\����_YSVC@ΤI밷7���s�ҕ�*�+N�AZVV��:df�j�1V�8B�^>L�ҭZ��@��矛����=�����B���3���,Y2��#W�s�Y��)u��v�65�cǖt��R�M*-����R^�}�.������7�f��;*E���#66���%T���&��!��)�P�+t��u��@GG���11�e�*䑟_yS�GEʗ�67/]T���E��d5��BEe���#9|8''K�N}�ѣ;�i^�D"������	ڄ�,4l����������!"��h����ŃI��2w�n�v���V4�,���.��;:�Wn��M���G^��O)+���4U
E��#nn�D�Y��	���beդ�d�iӺ�����Hd��I���N6*((,Wj;##�\ф�ܢ۷�jȚ������%��q��9���73{Ԕ5==�\W��BE�����,\���?���Ϸc��n���"����⭡]64{��K��ؽ�<����C���(P)�w�g֬�ޞ�?!b��)�\�
���Z�h�?L_4� =�W���ʕ��ƍd
e4ib����2���	oo{QeC ����̘���{�O>���U:~^��\x\z��rEʆ�=*Đ�&e).���/U"y���H�E�m낟�>��B&���T]��⾡����G��.ϲe���_��1c��6,�⼸�Y]5�m?	m)ͼf�q����k��᭷���ڣ9���bbb��e�:t6�bҤ��6Ic��0�kW/�v�Rn��/$22�+W�<��$�}�Yrr�������??G||���w���A��	O��ڔ-[��嗿���g�Y��y��02���H�V��
JO(����[�W��)�]�˅`m=�ڶ�<�WtQV��侲p���}�۪s!X��c�KU�TgNA��H$鑗WHJJ&k֜`Ŋ#��5c�����[3��U�uRv_u�����v�Vv�����m@.��h�~V�<ʂØ<���Mj4h��h�΍�^���x�/��m�mR���POٸ��LNt�=�\�W��5k����	@��Mzq"���[��&�@WW���HP�+�����W�Y�zb��V�?���ݵkO<q	���"���XX�9t�zMw�U�ye��yM���
���YS{��\P{�R�W1:�_}u��??���##Gv`���ښ�j�ڮ��~�*%�XEk�:��WѱڌTZDh�O��Ɗ�2$P�&5*4Z� ̚՗�G#y��-���p�Ctt$�lٜ�-�3dH[���������H�رH֬9�TZ���.^^v��9����fmm��w"���`?~���M�@��KX�<��=��m��ή�٩TZ���>]�zҧ�={z��l�֭[���{*�C�I���8UW��G\@�-�^���>�h���B�-1�)
%��U���uR�cR[7gM׻6��Aӧo�̙[l�2�T�@5h������o�ѯ�b�.=țoP�IZ���)ݺyѭۣhq5�����9r$�{����5���__G�����FT�hnn�ط�u�yg;�ǯf��~̞ݷA�(nTZ��ZT$�eK����Go:vl٠n*5�x��٣N[MLpp����66O���dre1����?�����3wk=}��X7���0~����c����"A��x1��a�ܹ�����M�^��k�n�����Ԟ�����,""���8|8�ի�){�(�8�aj
�S���AC��H��K������n.\��o�aiYqe4uR�ZZ�^>�����4T��YUKJ׷��Ϗaժ�uΆ̱c���}���T��r���	GW��k��׉ȵR=������F*-bϞ�T�c%(O�3 'v�С����������bc��Vt��J�M*-"22���D���	O�?��������R7�f����Q1a��81m���]���!�zG5��u9}�}-�����G���۔�^�e0xp�'�%�ĤV�O"���+��HN@�3#F<����4kf��f�JԽN���>g��b���qu�f����@R�hČD"aɒ1���9����/F��$A��ץuk'Z�v�dO����Ë���9p�2+V��P����Z)�8��j>>�uڨO �kڶu���PBC�1|��̚̬Y}�p����ec��Sѩ*cTe��\�=i���SQ�CI{�3�@u煹��0b�ST'^ɚ�����T��7������������ߚ�K�`d��n�=�F� �ښ��g#�>}}���n�����;;sz��Qn+.�USؿ�" pr����A)t���iٲ�F�Eh'��M����l�x�y�~����,_�����M�w'Rj;��Ư�8U����k2�����r��
����B)`���U>WU�U�O	�U�*۴��L&�O~eŊ#̞ݗ��~.g��Ҩ���Am9�=s�l�С7i�\������O#<<���D�^M��?��r�Q
eʊj>>�x{+JF{{�cgWq�Y��!��]�ر%/�����/Y�x4�V�Y�V���L�Ѕ�C�
r��J���eƌ͜<y�+��쳢�r}������ѷ��V�l�.��� GGK-Ky��"�]K"22���D��X������Y����Z�+xyي|+A���۞�~�ͼy{�2�{&Lx�y󆊰�
��0�ǝ?��γ61lXÆ��� �p�r�Z�&�����_~y���VA��(�LӦF|��x�[ƪU�y��6I���u��w��߱��������L ""���~��_<(@GG���5>>���8(=9���*oA�=��g#�޽���8s�6+V�Wy���SWe�bO���f���x���o�D�6άZ��衧&��
reΜ�|��~�t�x�\.(r�t�K�6�LNll*��
�s�Z"�w�'&�2�cc�8�
�    IDAT�lK{��SP�@�6�̘�~żyC�0�iu�%Z�TZ���g���L��|0D��S#�V� ̘ћ�����7���"|HP)::�ܚ��֌���ss��J&<<���D"#�8x�
��+�F7o�|}�i�J�����аQ�j��ђ;f�t�A�'ǏG�x�hыI ���4^zi#��I,_�h�5�F}ť�#aٲq���s��⫯ƨ�$��allPa����,"#ծ]K�ԩ|��I


����ͭ���@񏋋u���.���t�3�?]�z2s����K���kW/u�&����0{�O�ښq��xxب�$�\� �ښ�t�&N\G��:T(hA�)n���3��ʸ}�.����l�v������Bռ��E���U�էS'w��sＳ�Q�V2iRW����6M �|��~֬9��q�X��9�рЊ�Dp�'v�w�Ӯ�[�4���t�����Ӗ!Cu����'**���eu�#G"�{7PTU��U+;�������[4 <K�&�Z��v����wq�h$˖�#(�UݦU�����m����E�l߾��C������v-�W^�̝;�Y�l�=�N�&	� �kI����B\���!�w�*�j�������Jz�4���$��� pp��U+;ePoo{��#����BC⯿�x�^���o0�bϜ9Cǎ�m��1����n34��s�h�"u��6tt���z���s��^������_:t�P�U�\�ڵ'����8�l�8\\��m��<3�F� DE%1`�WL�ޝ���ns�
���ϵkI\�����ZQQIH�E�����j�����2\�ͭ�(-@.��i�i,؋�[3�.[�4�@ ����p�>~���[;��Cx�i�'��������o�n����9��8�6\�K� l�t����ɶm/k�L����7 �v-���bcS����)�q����pr�T��5}�7����go��+�x�~��@ ���X�hG�F2`@k�~{ ^^v�6���r�l����bccƲe!�	f�G��������<8��͛�������I��JR��)�֒ILL��̈V�Joo;�G���l�p�O>ُ��K���]���K#'G�F�h�>���	�Lhh�{����ǜ9�8s�/�ؓ��~��,���N1���G���qr���_�CA�##�2D-""�a�D22 `mm������x{;<|��Ҳ��-��������vN���ԩ����E�3�@Po�dr~���}����̜ٛ_��`�Ba��5k���pw�aɒѢѺf��b�ʕx^ʌ��3����ꅤ������(~�_O"3SQt�y�je��������ssєQ�������̛�c>�d8=zx��,�@�E���z�q�/?���	���9��Z���>}����It�=^=�3z7��)�*��b`��Ӽ��N�l�^�_�@�m$$�s���{s�z2׮)�ֲ�Սlm��	//;Q>Z�HN���v��E�i���ð�5S�Y�@�HN�䫯�`�������Э[�6�MN�d��=��F�^�,X�nn������n1��+�9y2�?��#�
e�s'��Ix(r��~=���ȱ�3�U��"�OO[�65R���q�P8s��"=�o�=�^�ֻ��@���Jb���>AϞ�|��u^$ /O���'Y����M�裡���_�s
�!f���0`	͚��c��?#<�\Ν;iʒя�Ւ��- ���RY]M��c���-���j�^PLnnK�d��c��9��g#D��@ �wN����y������y��*��dr�o��/�����^~�'3f�n0y;�Z!�@DD�}͔)�x�A�6G �Hd2��9�DE%+{�ܸ�B^��D���B�je�[�����D$�����D�yg��E3~|g�����(!��L��������HO�K/�䥗zФI�o�>��E��q#�ѣ;�_��6.��)���aΜ�ٴi�{������PT$#.�>�����r�_O����D���^^%���e'���>��Wrs�����	錞��T��#/O����Y��������@F�h_���#G"X��OΞ�̀�y��Axx�ԁ�5#�LI^}+��s�`(���٠@P�Ɉ�I-'rn�HF*-BGG����R���xz�bh(@�99�,Y�kמ�E��|��󢹰@ �w�����/��Ӳ�~�,={>��\.����|��A.]��W/�x�AA��V#F�����0`�W4mjĮ]3Ey>�@ʈ��ǵk�ʼ���dn�LA*-BWWgg+||����U������]>���y�A���;���~�}�.�����<�L+�����c��


��0V�>FDD"���3kV0�j�ZP�1S��ד0`	��uf����6G <D*-���Ndd"�oߥ�P�������[�'���F��r�h$����֭F�����}��Z �;��s�E���ȑ퇣�%IIl�t�~8MFF.��a��>��ث�dA�!�LE���K/mb���{�����A*-�ƍ�_O"22IYJ:66��B�����=9�ak-Z4"�
�drv�8��ſ����/t�ׂE� �@P���r��	��O#))77kn߾���	!!O3~��"�_;b�2���æM�ٻ�5��ʻ4Aæ���7R��J*��w��"��qw����OO[��l�������S���͛O����w�q9���������(D,%��F���߰9�6��6c3;o_���f�洍09�1�,�$)*:����԰RRק��~�uK��9<�nn}>�����N���fҤ��6u���֭���
!*��,�6���_�ιs�03Scmm��V�LXRiI1S�����.�ʕ$v영��<��"���q�B|�9��9�H������so�#���L��׿�d�^45&��|�o��}���0!��� �s
!Iddk�a��#��eѯ_sƍ뀧�_~����è[וٳ{ӳg��
ӓb�a����S�����eAM!*0�V�ŋ	y�FGD�̬�@v��Y�˫�}SHׯ_�*UlNoz�ne�t�^V�܏�``�h&L�H��U�v�mڼ�^oD�VѻwS-)-_B��JI���O�n�Q���fM'��c�ȶ���߷mT�M���Ɩ-Ѷ���f�_�H1S�S�b8�KƏ�Ȝ9����M�:9��qDF�9�SHgddP��=��nw����Z5�B�^���f�������IN�`Ȑ�x��ԭ����`ѢP�Z= ffjZ��dժ� B�`0r��֭;��� �ݻ)Æ��߿~���ǏG������+Ђ9s�ʄ%��3E�n�Q^zi-K���o�fJ�B�F���W���L�뮖[�ܾ�@�*6�uS���)xj�rB��Xݭ��u�_�ŋws�J"�z5���$'gܷ�Fc���k�>O��
�B�QQ7Y��!!ǈ�M�U+O�kM��-pp�z����q�������oԞiӺ�VTR�՜9?r��[����t!D���JD�����MD���
���^^9]�r��y{����\��Y?�p+��&O�\����2�l���JD�u�����húu�Ӡ�L�*Dew�m�N�u�_;v�j�x��'6�5^^����V����p�o ��RF�j'3XVLR��V�g������ʎ/�i��r�};��:9�y�DF&����/�jxyU��S�~�[+�F� 89�0sfoF��+������8v�2z�!��55�Z���^��AQv���b�ֿز�/��3
;;+z�lL�~-��ɧT䤤����w�r�~�ܪ0wnz��I*)fō����)��`ժ�*\7!�2�Ҳ�릖[��N#�Ѩ�]��n7�
/����X��޳��ӥ�FG���G�~�K��Ydd�(��V�P��,Z4���[����eõk9�֭q�x���٘>}��c�����d>�`+�7��e�ڼ�� Z��c�s�R'�̣:~<����������=��#���r��y�йx1�V�J��V���r���ݝ����Z�O��B���{M�Va4iذo�5����H�7��ȪU��?Ln��[�81�D�/�P΅���y�;N��W�
��}�ӱ���]�N����w�С���׌ٳ���YU�<�DH1S����93�+�ѣGc��!*��@t�MΟ��o���23� ��U�g�7�]KfѢP���73S����ћ7��O�Ə�Ppnw63��
/j ��o���7Z֢����q��BC�ٵ�,11IT�jG�n��ӧ):([���_N3o�v._��������z��3���k	9�֭�����t!��`0�t�x������l��.,����tFh�k��!..�6m�<r++o�͝Q�,P�,P�-Q�,�~�@�� ,P�5���Kr��df^z�s������,�c�R�Lhh8���ؿ���Z�5�K_�vmHӦe���Ng���`�/h�z�O�����\�%
%�Lq�t�_�ŋ7ضm:nnU
�I!2b�R~��<�����G�1�h4Ү�+6��ڵ�J-�Vk 3SOV���L=5jؔ�� ����`6m�T�X)Q�ddds��e��"س'���8������]ҹ�o�]W+==�E�BY�t/ժ90{voh!��)fGJJ&}�.������_�ںhq���Z�~��W����k�HTz����1B��
 +K���Q8p�"9q"��@�n�ХKCڴ�W�Z1bc�Y��WBB�ҢEm��釟�J���b�qEEݤ_��i�΋%KFK%/�(s�Z=���D���Ͻ��Z��ш����u�ҬYmRS�����'�3�V����+���C�"9v�2YY:���Ѿ}}ڶ��߿>��\ə3����τ�EЫW���/��mS5J'(�<=��t��}v	��m���(I!�s�bz��J�F�Λe��َF�jФI-6����;^^���j�%�!JArr:ǏGs�xǎ]���+dddS������g���_�����jr��dݺ�ٳ�<Ｓ����ȑmy�^���+���)��y���Ø1c>>n�J�HB��Z5����ׯ9͚y���NÆ5��,D%`0����D�����(.]����7�z�.C����ߋ�5���[ft�܀�ٰ���o租�dʔ.L��������=��)!C�>Edd<3f��NZ��T:�B ��lKt�'J�B�2��Htt"g��r�T�ÉѤ�e��hÓOz2xp+�z�.-Z����R��e�F��g�Я_s�,��_���2{voj%���R̔��^�Å���-[�IK!���T*U�cC��%E�7p�b�O_�̙ؼ�))w077�~��4kV�A�ZҪ�'^^�d\o1��Z���=9�-��ogƌ5,]����H�v^Jǫ�d�v�N6~�N�g����
�B��}@�REEe-f�����,11���8.\����8{6�s��s'kk|}�iҤ�פI�Z��֨P3��5�y����s��@_��폷��ұ*+� ��Y[[������s�~�}733�ұ�BQ�%'��W�DD�s�|II� ���Ѡ�-[z2fL{7���Wu4��0%oo7V��DXX��3]�~���~̘ѣRN��4)fJ���#+V�c��E���O���O+I!L�ޮ,>�/��֌���{����!�}�V�q
ʙ�q�;fq>��dz�ex���a��x|���DE����w�� *�&��	$&���dK�nԯ_��}�S�~u4p���N���^:x��//r�~���3uj '�ڃ&$�L)i�̃�����+�YӉ�S��$���a�GaE�ö}T�ZŃ�z/�m��'�s�w�G��:�(:��@||
W�&q�j2W�$u�K�nu��7s
ss3j�r�nݪ4jT����S��>>n���+�[��R�U<�Ll�ҥ{Y�(�o��ϬY�:��L`R̔�������y��qq���g���$�&�(7�m{oab��G=��-���a?��8�IJJ&�񷉍M��u��W���I"66���o������vm�֭J�9���֭��gUj�r��a���9Ӧuc�ȶ,X����7��cΜ~t��@�x�3�l�Rx������ѽ{c�#	!�0!�g�R���V�'))���t�_�͍����&!!�{||
		)�ǧ����������5��U˙�kҭ[#j�r���ժ9��_ɸ����O3vl{���ΈK�ܹo��_�Jǫ���1��3{���������/вe�#	!�0�[;�>�)i�zRS3II�CJ�n������IRR:7o����q�pI#))��7SIMͼ�8VV渹U�Z5�Ww�iS�Ww�Z5�U��ͭ
5j8Ɍ��@��n�X1��#y｟����mͬY��$ 99GG)��H�y������f��%l��"���JGB�RW�q R��Yi�[�q(�<V����l ���dd���`0�W<ܾ}'��))w0r�f����ΝlRR2��Ғ����zFF6ii���e�-^2�s';�,���8;�R���ζ89�R�nU���pq����''[��mqs����)�d�k����3ؼ�|��͛O0qb S�bk��EKϟ��K��<���T q�#Ō����Y�d4�G�ȑ�غu��J�B�����{o��ރ����7��6N�q>���Vڅ��ujԘQ"ǲ����R���%vvVXYi������kk\]��y���{���9_9��R%�uY"A(I�R1p`Kz�l·���~c��#̘у����;��ۛ ظ�8��RE �f�XJJ&�}@H�2͢��2�"�E�nY.YeWpp0�GOf��} XXh��ə�V�Vco��Z�R��`�����UތO��V2(^TxII�,\��}w��u]�;�?�����E0l�Wy۩T*��{�Q��)��̛*Ō��n1p����ڳ~�2��L�bF<
S��"����{��̎�i�֋��[��$���Q�U�X1N&�*�Ty�� wwG֭{���D������
!���J�ʷ��}=����q�SR�Z!D��������زe:ׯ�&:���	�F�8q��PʲO��xzVeժ��`ƌ5�$KQ�=�o��h�������z�s��qJJY�#�(]��kF�\F�����K���i�d�3
jٲ˗�y�	���q�B!��-[�;������`0���͐!�#11ʹ��)f֩S>�|8˖��'���t!�Ba"7n���g�:�@���K�����b�8�%<��cѢP��!�Bػ�<YY:4��Y�
���9w.�Q�����M���ufʈg�iCf��9s~��RÄ	JGB!���w�X[[���q���q��Ubc��덨�*43�Z}ޘ9�NϡC��6-�ŋG�� H1S���OV����ތ����+.�(��t�
E�U��Q�L7��h��[��2��(�'��ׯ/��
Q���Zҷo3�|�:3f��vm=*224dd�����ݜ�l3�ƜI6m����РA�ҿ��xyy����u)fʘI�:q�N6�go��Bða���$����t��3�<�^/�JRx�ffF4H���4S�gfj�x�
�#���8;g�䔉�}6%�`wȐ!xyy�����dv���ڵk2d*�[[-��Z\]��F�Wq�NN���hM�j�6�܇%R̔ӧwG�3���k1<���ґ�����k֬Q:F���_1��5�ny��qww4�y��t8p�]��ΩSI����K``C��`e�,B�����(�L�]�7?R̔Q����
^y%���ȑm��$��4k��֭35j�{�?L�Q���~^KK]��ҥ�/ ��q���c׮s������*ڴ�G``C�woDݺ��Q!�'�L���=13S3k�zt:c��+I!D	�Uˉ͛���s+8�K�,C`��I3�������ԩ�ܺ�������y��?��;�l�n]W�ukH׮�hӦ��f&�'�E!�L7}zw43�������q��$��88X�z�D^}5��c������c�  IDAT3f�2�m<���B�3���ٵ+��fٲ�qp��cGҵkC\\��)��b��:5�Z�ܹ�����󝕎$������p�ԩ����Ht�M�x���M�&�F�����=�o��ʕDBC���og�={=Z����kӵkN�M�F5dzX!�b��)'^x����|s7n�0wn�x!D1}zw�ԩʌk�r%�E�Fbee�t, j�v!(�AAHO�",,�]�αj�>�h���ҵkC:t����B��B�"R�Tyk�<����9���H1S���;�M&!!����>�BQA�w�*������b�8�ܪ(�>�����ل�=�`49}�j^w���Ø����_��]苇��ґ�(��)H~��X%IeT:�xd��G0n�
Z���o����T:�B�r��Ǝ]NJ���f�Z�Q:R�$$��{�9BC�ٻ�<��Y���獳i��33��1�(�r�6�m��HAɽ�e�����g�3�ԙ3���77G��~���JGBQBRS3�2�{��`��!�ne�VϡC�y�6QQ7qt��K_�ukD@���6J���(n1���+�+؃EJ�{���^+�b&����H1SAEG'2b�R�zk�L�ӳ�ґ�B���ȼy�X�x7�=ב7��_n[6"#ع�,�w��ȑK <�dݻ�4���M�B(�8�̃�\�V��ZS������3Xbb�F}MLL˖��m�'��$��m�|�3�кu=�,]�[4RR2ٻ7�]�αg�yӨ]�%o�N?�'���!��ry�b���K���OQ���&�L�����������zk@�k�FE��BQ<�O_%(h9��v|�i����<y��~;ˮ]�����%:xӵkCR����1�(u�Q�<��]ƊS�v�ߗnf�_�F#��2�v�y���`a����N��s�b����̔�B!��ƍT�{n%���X�xݺ5R:R���M&44��;�p�@$YY:�4����iSy('*��n�y�~�^�b���?j��<��)��oſ�T*��|��s��q�A������y���>.\��`0��{?+�T!Dq��ڳa���oAP�r��b��S����5�=��?��g���o�Ӽ�k��wl�/�����O����t\!ʌ��,�ڄ2%��4�F���
�ҥ�L�l�X��-���S�z��*8x>
'BQ+W���[��ݻ)<��mş����ػ�6g9q"335��y�uG�IpDyf����'��=��2��(1������jv���՞��t��bF�V��lþ}�����BQY8��ɫpr�aٲ�4h�t$�ILLc��pBCϱw�yRR2��F����ŗ֭��<Z�ӧ��v��M�N�j�܁0��Xg�,,`YZ��Y%dooŊ�x�z$$��2 ��[�����L(��q��{�s�+���ѧ�g�[wT�H&��bǐ!O�d�Μ�����ڵ!��z���^L��o0y�w���$%�阛6��ʕ������^ʿ���4�n�'R�T`[��šC��t�����ٶ�/~��ɄB�7�*�_?�q�:��Kky饵de锎eR�������{������=HNN祗�Ҭٛ���_~����kg��S@��ѣF}�ܹ�ή\��(_r���~U�V��H7�
���d:u�OffC�ۨT*ll,���YԨ�hڀB!J�Νg��V���̲ec�[�U�H�KK����ϳk�9v��ƍTj�t"0Зn����9QQ7i�����h�ԫ�ʲec+�Tآ�*�nf�����5�CrrF�ۙ���䓞l�0E�+����r%�I�Vq��>�d��5W:R�a09u*��;sִ9s&++sڷ���[֬9|_�l�)h�j5�;�ѣ�)�\TR�<����d#��9O��j�Y��j�z���7��3U<!���vm6o~���~�I�V1g�Oh���j\��*�7��̙���ח��Ϸx�A��*�̷�Ng@����k
ZNrr���!LG��
H�V�m�t��?`��Q���;;+ �%�A�����BD�uSGBQ�,,4|��`�.CH�Q����d�c�9իWa�p?-ITT"��d�F�F#�������H'B<�3X�*6Ђ��o4����OS�0! o.����ez��ɓ��'xBQA��ל;^"==����k�9�#�Iaa���_�t:=IIi�?�����.iBeȘ�r$&&�Ç�ȱn�����dN�J�ҥ���5k����J����J�B�b�s'��_����c<�|gf��o+}e����ذ�X���N++����E�Z�h۶��1�%wLHHH��Qʤ��`6m�$ �w�ƍc�ʕ%~\��K�:�����Ij��?GyĊ+��!��mݺ����OxyUc��Qԫ'��Ԩ1 �F�V�T�TE�r��j����N<��z[{��Qڴi�X�P�,�����u#,-=HN�Bf��J�<���|Y���dĈ �^�Z�$��|�B�����L��.���y�Y?�#)6�V����@H��,YD�*���Xbcc�����lg'-1eQe�,))��~;Ö-'	���`��ms���8;�*���M�(�@!��Q��+�7����`����9���J��)�w97�+W��ȑ峛��<��o�}�i�l9�ѣ����Ϲ�X�T*�.S
 ��B!*ss3^�/x���~�_��];/��	!
�ȶm�e�IN���Z��`0�m���5��܌n�ѷo��,ŌBQ	��{:�W^Y�С�c�� f�ꃥ��QV$$���o���h�����9��>H�Rakk�GU �rdjf!���rt��o����g	>L����c	!�JK˼;�
�.��y��>Vi���bF�;*�J�BQ���wϢZ5����O>�E�3!�J��׃۔ֱ�J֒>FEP��+˖��ޮd�177�W�&��{Y.)fD�S�f*BS�QÑu�&�����=���ו�U!�w�n4��u�v�^��F��c?�G�*_߾�?�#M���*�
kks��b�de�3B!� rn�ƍ���]�`a��G�,^*����)S���d[`A3�P�V�3q��A��
.�IIA���mr.�i�Q�W�~Ei�~��PM�BQ�ԭ�ʦM��Wz��'�Ч�BΞ�U:V�t�5�(ק��-�y���^�r}~Ԭ�,�y�?BC���s�j�?����ݻ7b��
&T�3��J�ʷ����ɹ���{��+�8E�R��O!����2%�]�fbmmA�^�2o�6��tJG+3v�*������X��Cɯ�V~�?��������xG��w�N6����ѣ��C���W_�Λ@���^V�f/{�3�����>���8NQ�/��pO<Q��~��;�bŊ0�v���G/)��y�kLI�k)n�d��:C�ظ�_}5�/����ݺ5���;`0�?(���
�U�3�XJ�{Zid���G��!D��*��ڳg�,��qa��E̙�#iiYJG+�Lu*�z�_��8Y�r���=�y+���g��F�~�������3�߿�}�̞�oo7���W��e�de,Q,%��Rv�����BO͚N���D~���|s;v��wү_��w��Ly�y��]if�͓_.�.�#<�ӧ��x���Ǆ	�-�45{��R a�$-3�=�`Ò��A�B!J���ߓ���F�N�<�;�}v	QQ7����®9�yM*�c+u����m�Vϧ��JϞ�beeή]3�81��~�J��J��f�>1�~�=fi�O!Dgg[>��6n�JBB
]�|Ă�V�	������{�a�z�u���{�+�����o=��~�>{6�޽�x�n�x�7��z�\��U�H1S�֜[����7���{�G��Q~���~B!��u�z���+��jo�,�C���������e2��<���u��q(�m_�s=����炎U��7wy�����_��{!��V���d���]E#ŌB!�F�f��N��7�F�j��K?~E��z&݀Dq���.]>b�ҽ��f6l���gU�c�[R̈ɯ�[fBQwwG��z,�WO��������^1g=�nR�Qܼ�Ƌ/�fذ��Wϕ�{g1~|Gi�yL2����c,��qt�܀�����̟���1kVo�m]�n��)
c0	>�l��ւ�˃�ٳ�ұ*i�B!D��h�����9��ՄW_�g�<�t4!L&<�~��o��gZ��ﳥ�)aR�!���8;���O�k�L\]�y��Ō��╎&D�IJJ���7У��F���2o�5 [[K��U8R�!���y{��z�$V��DT�M?bƌ5��&+M����Y�d/��}����裡l�<��k(�13B!�0�Ν��ƍ���_����1c��6��ζJ���BCÙ;�'�_�ͤI��:5PZbL@�!�B��Z�����I��o�?�/v|�ɓ;1iRg���P��y����s���[�~�Ԭ�t�JC��r��Ғ�+W�t�J#((H�BQa���Ԟa�Z�|�>/��ʕ��<�3c��cooe�,666��#��ʕD>��W~��8���l�0�v��U騌2�`���Ç��Q�������t!��n��`ɒ=�\��Z���x8:ڔ��u:?��3z����%JG�Z�h۶m������|��o�Ys�Z��y��Ԫ�M;^NL�bF!�e���,_���ah�:ƌiϤI��Z�N�h�KLL�/v���qq�c��n��F��R�3B!�(��ӳ�,Y����,F�lˤI��Q�Q�h��m1\�<[[^|��F����L�hB�!�B�u��Z���x�nn�L�O�f<�\GZ���t4Q�]���ҥ{Y��0���L�҅���X[[(M�C�!�B�Z��͛O��7�8u*�V��0aB �z5���Ĝ=��Żٺ�$nnU�8�Ç�ac#EL$ŌB!ʟc�.��7�ر����g�?��d�Q<aa,ZJXX����Я_sS�I1#�B��+66��+��z�a��u��ߜa�ZӦM=�fY*%%������9w�:x3eJ:v�Q:�()f�BQ�edd�a��ԩ<=�2d�Sކ�ի(O�1�q�ի���'Q�U��3�Q��JG�F�!�BT,��q�[w���c��fҩ�C���G��XX�z�խ[��#8�0�i�ԃ#�0�%�[�U�()f�BQ1eg����3��e�޿����w���ӌ���ˤ�@JJ&���ض�/v�:����A�Z1|�M��R:�x|R�!��⋏�͏?��Or�TU��УG#��iF@����T II����i�o?EXX ��ק����\�V�X��B!D��Ķm�ض�$�y;;K�vmH߾����[[K�#�G�������q�C�.bnnF�N�ӧ)ݺ5���Z鈢tH1#�B��+.�[�����8v�2ffjڴ�G�.�ڵ!^^Ք�(�q�V��_ ,,�}��&::;;K�tiH�>M	l(��TR�!�B $&��w�yv�<Ǿ}s�V��؈v힐.J
���q�X���MXX�O_�ys:t�cGoZ��qP��3B!����8�Ν�س'��g�aaa���t�s�ܰaY˦��F���ط/����9|�w�dS��+�t����}��LH1#�BQ���BCϱo_��G���Nժv�o�M@@Nq���t�r-.����tۿ�7n���b��}:v��cGj�rR:�([��B!�x���gcٷ�o�����Kde��򪆿}����ϯ�,�Y���$��đ#�8|�"/&`i��u�z�С�7��D���/Q )f�B!Gf��#G.��C��>}�΀�gUڴ�G۶^��գvm��*�`0q�Ç/q�hN�r��m,,4�hQ�6m���_�֭�ai)�d�"�bF!��$��g��Q9r�C�"9q�
��:�ܪвeZ��M��uhڴ��s�G\�-N��W8y2�S��������O=U�֭�ѦM=Z��-k���!ŌB!Di���q�D4ǎ]�{s���o�V���N��4k恏�;���89�*��t:QQ7	�FD�uΜ����+�ǧ`f��ۻ:͚զE�ڴj剏�ffj�c��C�!�BS�~�6'O^�k�8s�*�ne ��j���;>>n���Q��+θ�;��(Sܾ�Attb�WD�uΟ�#""��l�OϪ4lX#�xiҤ�,@*J�3B!�eA||J^��������8.\�'%% �F���#�xx8S����689���d���-�ζ8:Z�V�څ-##�VGFF6iiY$%����NBB
��i$%��+9�KJ� ��ͨYӉ'�p�A����]��n�ƋP�3B!�eYrr:11Iw����I���$��SHJJ#99�����777��&��$##�V��v�;��mqq���ՎZ���Sǅڵ]�]ۙ5�k"R�!�B�w��:���IN���-ii9�9Z��_����5j�
{{���NN�8:�(]��!ŌB!��\�*�B!�B�rI�!�B!D�$ŌB!��\�".� �t�    IEND�B`�