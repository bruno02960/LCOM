<map id="rtc_subscribe" name="rtc_subscribe">
<area shape="rect" id="node2" href="$group__devices.html#ga82cf81704efe26b2e078804bfb67f924" title="devices_subscriptions" alt="" coords="153,5,303,32"/>
<area shape="rect" id="node3" href="$group__spaceinvaders.html#ga3c04138a5bfe5d72780bb7e82a18e627" title="main" alt="" coords="351,5,401,32"/>
</map>
