<map id="rtc_unsubscribe" name="rtc_unsubscribe">
<area shape="rect" id="node2" href="$group__devices.html#ga916e9be5016bede8624ac7c89f9eda8b" title="devices_unsubscriptions" alt="" coords="168,5,331,32"/>
<area shape="rect" id="node3" href="$group__spaceinvaders.html#ga3c04138a5bfe5d72780bb7e82a18e627" title="main" alt="" coords="379,5,429,32"/>
</map>
