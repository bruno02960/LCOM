<map id="init" name="init">
<area shape="rect" id="node2" href="$group__video__gr.html#gafa847549e9dc6e4f49f651623bc456dc" title="Clears the buffer. " alt="" coords="822,144,910,171"/>
<area shape="rect" id="node6" href="$group__xpm.html#gab41dd197773f68e69e18c73a8119ba5e" title="object_creator" alt="" coords="472,588,576,615"/>
<area shape="rect" id="node9" href="$group__mouse.html#gadd35ac18db20624e86b0c104a02fbf0d" title="Unsubscribes Mouse interrupts. " alt="" coords="92,524,231,551"/>
<area shape="rect" id="node10" href="$group__game.html#ga671b58f5509a3a9fa692bacccfc32cc9" title="Receives drivers interruptions. " alt="" coords="118,473,205,500"/>
<area shape="rect" id="node16" href="$group__video__gr.html#gabdd05df698103c4641478f491e11e284" title="Copies buffer to video_mem. " alt="" coords="796,245,936,272"/>
<area shape="rect" id="node26" href="$group__mouse.html#ga7528b123a3779d689c06876b78a0b91b" title="Subscribes and enables Mouse interruptss. " alt="" coords="99,575,223,601"/>
<area shape="rect" id="node27" href="$group__mouse.html#ga91fe374b9624fe2a223be3af605b1dd4" title="Sends a command to the mouse. " alt="" coords="99,625,224,652"/>
<area shape="rect" id="node28" href="$group__print.html#ga5f04c1438b5689bedddc17eb0dd9d060" title="print_message" alt="" coords="641,144,748,171"/>
<area shape="rect" id="node29" href="$group__print.html#gabbb46faef7390f85ad76868944abcf20" title="print_score" alt="" coords="481,245,567,272"/>
<area shape="rect" id="node30" href="$group__file__handler.html#ga90d3bc0149cb0d2782d63aa42cf3fa86" title="write_score" alt="" coords="117,1005,205,1032"/>
<area shape="rect" id="node3" href="$group__video__gr.html#gaa55320d571dc2cb8179422a9d8114de0" title="Returns horizontal resolution. " alt="" coords="1144,448,1216,475"/>
<area shape="rect" id="node4" href="$group__video__gr.html#ga36218c155eade74951ce7ffd60711a9e" title="Returns vertical resolution. " alt="" coords="1144,296,1216,323"/>
<area shape="rect" id="node5" href="$group__video__gr.html#ga5c30cdd3eab0edd2734ab3871f7000c7" title="Returns number of bits per pixel. " alt="" coords="984,245,1096,272"/>
<area shape="rect" id="node7" href="$group__video__gr.html#ga1cd7727ad0fc3fe3ffbbb98cd9115c1c" title="Returns a pointer to Buffer. " alt="" coords="1003,549,1077,576"/>
<area shape="rect" id="node8" href="$group__xpm.html#ga05b2c5e4dbcaffa701703b50a2111783" title="read_xpm" alt="" coords="1001,397,1079,424"/>
<area shape="rect" id="node11" href="$group__xpm.html#gac0e395e7e8c65b90f0680c7a917f1acc" title="title_creator" alt="" coords="821,397,911,424"/>
<area shape="rect" id="node12" href="$group__game.html#gaff72f275b5af37960b3baee51f855041" title="Makes a game round, where updating action on screen. " alt="" coords="315,347,370,373"/>
<area shape="rect" id="node15" href="$group__xpm.html#ga8b990eb150243edd20fb9c4182748528" title="buffer_destructor" alt="" coords="807,549,925,576"/>
<area shape="rect" id="node19" href="$group__game.html#ga425ea598437d36368c0e136f2be75a61" title="Makes enemies down movement. " alt="" coords="279,701,407,728"/>
<area shape="rect" id="node21" href="$group__keyboard.html#ga6d2cc119f3d1b28fd79e7acf2f4d4596" title="Reads scancodes via KBD interrupts. " alt="" coords="303,448,382,475"/>
<area shape="rect" id="node22" href="$group__mouse.html#gad34fbf075c41898c2120ed2d0ee6b20f" title="Reads packets from mouse. " alt="" coords="295,499,391,525"/>
<area shape="rect" id="node23" href="$group__mouse.html#gaab4aa4fb914d5e1046d1391b97091546" title="Checks if the given byte is a mouse byte. " alt="" coords="287,651,398,677"/>
<area shape="rect" id="node24" href="$group__utilities.html#ga88386f4f23c71aba0d4e995a5246f981" title="Converts a number to its twos complement. " alt="" coords="279,752,406,779"/>
<area shape="rect" id="node25" href="$group__game.html#ga1fd9e64dab3abe9facfb4dd7e1267bae" title="Creates the pong and switches game state. " alt="" coords="305,600,380,627"/>
<area shape="rect" id="node13" href="$group__print.html#ga1243268c621c2049a41956ccfc934fd5" title="print_info" alt="" coords="487,347,561,373"/>
<area shape="rect" id="node17" href="$group__game.html#ga9a691a2142903ae9009a88a62464ddd9" title="Says if there are still enemies. " alt="" coords="478,397,570,424"/>
<area shape="rect" id="node18" href="$group__game.html#ga8aead8655bcc62fb760afdf2fe161ab0" title="Destroys the enemy hit by the pong and desactivates it. " alt="" coords="655,549,734,576"/>
<area shape="rect" id="node14" href="$group__print.html#ga4316256507429b01e848fd72e5fdca73" title="print_number" alt="" coords="646,347,743,373"/>
<area shape="rect" id="node20" href="$group__game.html#gab806d0bb50ec52aaa6ad9a71a2d3a05f" title="Says if there&#39;s an enemy going under the ship. " alt="" coords="493,701,555,728"/>
<area shape="rect" id="node31" href="$group__rtc.html#gab7e8ff751e63b72d14aa5f7ec727d337" title="Returns the day on the Real&#45;Time Clock. " alt="" coords="311,904,374,931"/>
<area shape="rect" id="node34" href="$group__rtc.html#gad751c36263a847ec77044899618cfd66" title="Returns the month on the Real&#45;Time Clock. " alt="" coords="305,955,381,981"/>
<area shape="rect" id="node35" href="$group__rtc.html#ga37f344d06f4e1b826aed5adf7b729fe8" title="Returns the year on the Real&#45;Time Clock. " alt="" coords="309,1005,376,1032"/>
<area shape="rect" id="node36" href="$group__rtc.html#ga57e0eac5ae1c791f2c63b0740ab94e08" title="Returns the seconds on the Real&#45;Time Clock. " alt="" coords="311,1056,374,1083"/>
<area shape="rect" id="node37" href="$group__rtc.html#ga59e635249f9555c53ddc24e54b82f01f" title="Returns the minutes on the Real&#45;Time Clock. " alt="" coords="312,1107,373,1133"/>
<area shape="rect" id="node38" href="$group__rtc.html#gaa14f12da2be63f2a594cadff28d10f40" title="Returns the hour on the Real&#45;Time Clock. " alt="" coords="309,1157,376,1184"/>
<area shape="rect" id="node32" href="$group__rtc.html#ga0eacd2fb5986b142e032ab0f8365a542" title="Reads content on register. " alt="" coords="488,1005,560,1032"/>
<area shape="rect" id="node33" href="$group__utilities.html#gaa62d5f8252ae370122486e82d3fb7de9" title="Converts a BCD number to Binary. " alt="" coords="455,1056,593,1083"/>
</map>
