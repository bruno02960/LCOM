�PNG

   IHDR  �   =   ؘ�   bKGD � � �����  `IDATx���{t�����			����kC"`��(��DKZ��h�����U����S�-�h��m)=*��AP�j B�H�!���n�����4	�����3��~������|3���of��QX,������/(E """""��'""""�#,��������Zt """[n�lBm�MM�0L����b����	 �j�jj��

���6�����Z��������7o�Ы���

@ppoܟm�\�������8q�EE�q��5��ע��W�Ԡ��٥i ""��}1rd���1c!,,H⿀ȶ�#��/ ?���W�ܹ*\�|F�١��Ã1th8�s&L��G`Р0�&_��]t��ț�zv�>���((����
&DE�aذp���GLL���Ghh ��zA�Q!8��j%���B�@}�f�z�z�uu:\�Z�k��Q]]���Z��^Eqq%�_o�B��m�E��b1y�HL����ޢ	���#���k�i8P�����z���؁��鏐��

@`���Ahn6B�oACC3�QVvee5�|����'ʠ�0z� ̞=�g�CLL?�.�|""�8�ɌJ��S��;OA�7`ܸ�?~X���C<�����9S���8x�EE��V�����c��	�:5�ʣȿ544c��شi?jk�0c�<��hL�>���nO�`0���v�8����~�?��O��_��ȑ��/X����f���ڵ�PYY����9s�#9����Gh���f|��	dfáC���^����{X��v�.�ҥ��Nׂ��ï~5ͣ�&�۷aݺ�PZz�'b��$��5��'""پ�k�|���<���x����NP^~���Ejj>�[o=��3o�|��`�oda˖|̝;o�9��޻��l�`��cժm��鏏?��l�3��DD$���f��jv�8�G�e˒0th��X���Ś5_`��#�?"�z���d�d2cɒ-ؿ���(fͺCX�+Wn��g?Buu�ҞCl�@aYH<�DD$��W둒�55�X�.�'ǉ��]�Nc��tDG�ÿ���W�Ȓ�X�<��Ǒ��<Ǝ,:��h��r�v�\��}yyO����$QW�ǜ9�P(��'�Bdd��Hn)/�������� �����S'۷ǋ/�"#c	�k��8�t�̚�F����O��C��I�DD$��_���Fl����� ���/����V刎C2R_�ǪU۰xq���{ ��M��s�i��_�a�ODDn��)��_���MO#<<�0�{���ED�����u�8pNt����? �ł�_���B[91�GX��^�񏟉�B���'""�X,�Y��nTT��3�|���ظq��h�;v0�|�^���W���Ll�v�'����0o�z�*��睢cu��r��JK���B�f�DD�o�9���&l�~[��Z�z��d�y�{1mڟP\\�Q��D�!jj��W�/�8�����
�
Fc�/U��z�	;5*
C����/O!6��q��X���jk���}�|r��P�U0[�)�&h4j����N\\$�Ãq�p)�f߾o��K��~�
�T*ۻ��u���K�<�$fW���g+D� X��S���4-� J�����⾍����ﻊ��DII���e~��k�  `6����d� ,L~�R<�?���D� �������o]������z��x�F���Ŕ�y7>��������Ʉ�}���1��/��{,����)>x;6n|���b6[������^>ն���K��m�&����;k�D,����i�f݁e�fv�ӑ�3���h4���
�GG��B$$���W�l�w �|��K�1l� �1H �DD�W^y?��P�UV��t��E���K���cʔ���� /�� �l�;��dbD� X��K
�{�q�i�rs���iiG0q�DE���B��TJ��~h뷞ɗ�E��O����S�ĉ�B��'""�࣏~���>P�:�R��Y�%�����8�%K��6l �zkN�����"ۜ�B���؁��� ,����-QQaؼ��P��Pt�|���Ί�����G��B2�����x4��v��ӧ�����V_�Gj�a<��x�QH�DD�;��u����?�Rr��#س���X���������&���-8Qg|p  �䓓'!QX��$~��;�t郲:����KX�2�'�'?":����!X��qX~�&��9���ذa/�}v*BB�u�A�����$�t�L<��X @qq��4������O�����7�yHt����̛w ��r�bE��C�xq��($��ҥUVUU�W^����?�Ja��HNN�%���زe��~���3T*֮]���H�Q\�r�J�����!�٬��C�  �'�N㚚�޸t)		סV��'����b��բc����ɤD~~M?��c�q<�g���!7���yq�'����<�lϞ=HKKôiӼ�M�����F�8--Z�����/i�Z�IKKCrr2RRRDGq��o� �\�ޠTZ0iRL&����=��k�B!�3�ަ�j�g��zƓ�Je�=�T�b�G�4�ʂ���=>������������z<�ܩT�f�KRRR���*:�_z�'����ɵ}��Ō���>{�B �~��_l����EG�;��.��s�����^!""""�[��'""""�#,�������|"""""?"�?1��=[m�O��D�c���&<��-[{�3ˢ�-7�<�)r��ڍ��k�w��[�KLL�޽{��ez���Ex��hll�k:>J�<�ZZ�ع�/ތ�7�D�q��s�v�����ƍ��z���K4G���$�����?���͇DG�8���3�-8x�K�lAI����䭇�ټM&9�h4�oJ��}�}v:� �h�dL�8Bp:�d2�СRdeCn�	45��͝;ӧ��η������'��^�#G.�ln�h�\9Kp2������}�qdd�ɓ����
NF�]FNN!22���� 0j� ����C}�d~ۙ����Ϻw<+��~�{]?�q|[g�M��a�M����}�م�yS�F����v�P(n9�j�����3G���seX׼�d�Na�%��"+�jj�Ѩ`0��ӡ�.��߻�e�u<w����u��ػ�[�ͭ�\[q��<DptYZk���sv�w7W�1[�l�v������|�نt�S�ejﵵ�殺:=���$22
��_
�R���>��؁���[�.����*rr
��~W��t����yeO����'wI��;��u�i{�j�mkz����Y����*DF�QTW�uj�C�zڡ�����{�:���:���
99Ǒ�~�]ڇ����[���6�,�ь�!;�>��$�z�ńoPw�j۴6�+��ځ��<�c�U�w��پ�RCR-SW�z����ؽ�,23����v:�n;��\�WQQ�m�Z���U����봧�'�����wu���}ޕ�^�S��
Z�Q|���~�h��Ř�3m��v6W���YG��J�_�[�����P�U0��}X��v���c�ʌ�_��je��5����h�j��;�vp&�t�bk����:�!s�;�Oo7=3}�����n�'���� �#���1ؼ�23PPp*�ۅ����nD�%m��[��w��7=)����gφ����Ѷop��Ξ���pUtt���E�pi��u��ɢ�U��j�G~~n�{mhw.���|�3��WE���o�)��߿���#��`0bРW<�aAAcEG�(��e���Wt���b����EJ�?;���vuu�,��^�����Q���Q������vxϱ��իw�!Bxx(Ǝ���y��ny����.8��g��+z��a� ���N��^�<	��n��]�6�:�6R�}��ϋ�L�O���4��W;�>^x�$$ĸ<o)�[�N���ij:�	�GU�7n49�lU*%���^Hhߜ9���Q�~��t7_do;)Ų��;���7p�Dt�f�T*��CC���ݞ�;������<�!Q�ZmƏ܀>}néS��gﻋ�P(0g�x$%�6���yt��������j�o{�ȅ��R*͈��Gj���ܹ*��B�=zK�jk�o��褥��kw)�Pw�j�R�>+�t�J������}�=����~ee5ݶ��G��NZ�|o�j4��������!/�<���aǎ��Z�R)a4Z��T*��|�����dr�̐�����xc;i0T#3s	ZZ�س�YY�ص�3
E{?��z��_����lntz<_m���=dHRS����&�o/�V{�O�w��5*Jx�HK3xm^���KR�w�wߵ���9[�ۛ����k�=��^{�����]�����.���8��7��Ü���F���-��e�f��ɲ�ۂ]�V���w<*�S��c��x�Y�(v�.Fff����}=m��c{���3�Z�ݙ��3c������4=řm����w�������444c��S��,@^�����˅�\��g���g�����!+�22
p��5h4jΟl�u]ېO���W����8�����7n(ƍ�U�~���:]3
���]Dbﵫ�9���aRf�g���;v0^�g����CV�1l�v͝.B�E��k[äZ�j<�Pz(�������� Z�kSS�$�ő6��w��|�}��x�f�nzRo{D,SOsGpp/̝;s�N@MM#rs[��?~*�F�UU����i\]3l� ,]:K��ę3���.DFF�^m��`K���R�F��wI�$[�/��*�S��a���q��������i�� QQa�ӑhJ��&���(Μ�=>��HJJ  .8�o	�y��BZ�s(*zo�9s�#����੧�Î/�ȑ7�b�O�V+1n�0��H�1c�����(,\�����r��_���$������xv��g��*_����F�3�`ƌ1������`,Z4�ME�伾y;�T��2%:���~<������VOl7J�w�=w�=o�=Wt��+]t�����+<�>�y}�v6��'�eJ����"�I���<��'""""�#,�������|"""""?b�"�}��y1�<�߿�>���n�j��={��~I��b޼y�c����s�Z-4��D.�j��#H�_�9��O�n)�ccc ����F��.:�ˆ����)r���9m�"_�����䈎B䖀� �\ֶ��6��q�'���
��DDDDD�7������ȏ��'""""�#,�������|"""""?��c�\N�i�    IEND�B`�