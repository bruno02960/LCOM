�PNG

   IHDR  y  #   �z�m   bKGD � � �����    IDATx���wXS��7	{�Ņ[w��Ҋ{/����[�{�n��Q7ZjAG�u֪�PDDv�������&��<����oB�}�9��R�T��������X�������H}򈈈���C�a�#"""""2 FB@�#((;w��AH$�^�vvvB�BDDDDT �ɣ�w���eb���8q��e{��#�����eh�H$�"""""�`O�a�#"""""2 yDDDDDD�!������Ȁp��	�&>Q*�TBDDDD���H"����ϪnCDDDDD��pM�YJ��K�C�H$�c����m���m�Җ�v����������pM*��C*U���-�N���P̬�GDDDDD�aO���Wv��<��Ꮘ���
3��F�{�$�ae�!�4J�=j��k��8\��&�Е�P�ݰˬ���PM""""*�ؓG��Z�O�<P�sf9�̩ZG/�������(CXN������}�|;��}��5�@؛FDDDD�[ؓG�ӐLm�<�������0cȣӅ`�5��$"""""2 yDDDDDD�!������Ȁ0�N�B���C��ݳܮP(�T�~,� �+!�*`f&�"""""�`ȣ�*U�T*E߾}Un�H��h�HM�����\]�)��ڐJ_!)���C.��U�V�ruDDDDD�'Rr�y�_߫�3g?��cÆ��^�N�r���7�⋅  �D�\��UK�S�z���:�_�<t'""""�Gي�K´i�
��ѣ[cƌN01ѯ����c�D���36�@*��xq+t��o���/�t���~=6""""�O1�Q�n݊��1^HM�a͚�hٲ��%�ۈ;���w!��?ۖ�033B�v5��7uо}-+f)@�DDDDDÐG*��q�_T����P����%HLLZ�\�wPd��O�	 /Ά�C	m�HDDDD�\B�>�w��7/ �'���{��< (^��V�6��\��D"FɒV([����#""""R��Q���0|�'S�q�4mZY��n�d��߀L���M �D077Ɖ�P�{񈈈�H��'�  �u�;��%�p���x ��O=Q��%��_��V�g�#""""�ŐW�)�J�Z��ݷ�[7g��;��6B��166fX�nTu`K$b�*e'��TFDDDD�y�XJ��G{a͚cX��7�/�cc��ei\��6�$��������P��:v\�B������(�xM^!���C����(���fͪ]�V%%��M�ex�"r�&&F�����P�'���?oc��^ps�B�R������=y�Px�t�/_�"0pb�x `nn��d,��paOT�n33cl�4'�Ǵi~�;�?�6DDDDD��=y�̝;�1h�f�.m��;G��w��}�Y<|�
K���l[``0<<v�y�ؼy(,-M������(o�
���p�NN���t��CKN���1l�6�+W^^#Q����%e�!���r�1ފ�M+c���055�$���7 v�.�@DDDD������=���Ѳe5xz�3��QŊ%8	66���m��}.tIDDDDDYb�3pǏ�Ð!�СCl�<�P,��	�JYc��	�V�z�X�s�]�Jy�ȑ�pw�D���v�$������ޣѾ}m��m���B�DDDDD���3P����8��-��H$tI��X�_�R��1~�N��&aȐ�B�EDDDD��!� ��s���F�9]��L$a���(^�3f�E||2Əo'tYDDDDD ����y̜��&��?t��6y����0g�?bc1sfg�K"""""b�3$۶���y�>�#&Nl/t9���{K�ؘ��c��94�����ǐg v�8�y�0gNW��F�r
�޽���c�z!>>�W�$7DDDD$.�n �칂)Svc֬μ6L@�O߇��v�jU[��rDDDD$�<=�o���'����;]N�w���M�T���;�iC�����3�#F��ܹ�ru�+W��iӦ�̰��� %%%׷ǀѨQ%l����&""""�a��S�N���C�a��fX�8��}�����������0���    y}�ܺ�~�6�aCl�>��zDDDD�<��C.�bĈ�ٳa�^f}���@e�G*�"   ���W�<|}ǡ_�M>�;v0��vp
@=s��S�..��re?NׯÜ�҂^pp8��Dr�T蒈����`��#w�<���&4o�u�q�~=P��=|}���ʹ����*tIDDDDd���Ŀ��Ā���쀭[9=�>Iz��Æ1��f1�遰�h�	���ؾ����:u���w��}��C�1���0��7o�1p�f�+W^^#ann"tI��������P��Y�]�|}��޽�<x+�iC���O�С�  ^^#amm&pEy�*`e���t)ԩR�VY�������4h��C���J�pw��ӧo��3%JX	]�I͚e��7D��m􈈈�H}�t�R����.��D��w<*V,)tI�D�d����o����n�T*U�_�b����sӦ��
�F�2ػwBC��涙=zDDDD�6y:hɒC
��m��Q�f���a��O���6U�-�m��nNmfW���W���^a�PO��ʄ.����� C��ٰ�~��V��-�.�3�m��#s�[~������fM�V�����ѣ� �ʅ.������C�ٿ�:-:�쎞=
]N�e5��r�fͲ�����b�d��
�K"""""=Ɛ�#Ν{�]�0�F�h%t9y�yX�.����c��������G""""�7�<p�VF�܎.]�cƌNB��-u�u�>d�a�?-Z8b�����.������C���¢1h�8;;`��:9�1=��
e���ڞ�Ǔ�~����an�o_�����Y�\�����2���,..C�l��C	l��cc��%e)����6U�� ?��v�ݧ.�ڵ>��R1e�nXZ�bܸ�B�DDDDDz�!O R�#GnGBB*��ss�K��Uj_�~M����9s�aee����]�	�<�̜��nE  `ʔ)*t9��t}9>�pwo���1c�^XX��W�FB�DDDDDz�!O ����ݗ��9\';�;aL�삄����`ii��
]�8N��eG����%���=���u�.���̙�1dHs��ӧ�]�8�<-�q�)ƍۉ!C�c��B�Czd��ѣ�ݷ����B�CDDDD:�!OK^���ȑ;��U�paO��!=#�������W51t�Vܻ�R蒈���HG1�iA\\2ڂb�,�~�`H$|�)�$1~�u0���cР-x����%���+&�+0i�7޼�Ǒ#S`cc&tI ��}����11f(^<Y��h�L&���氶N����<dl???����l��=֢O�
��%��.�����t�H�i5j�̽س�*��ƣA��Add$<<< ���|ߤ$#<|X�ߛ�~�hXZ�j�B�{���� �DJXX�`c�
+�TX[Kan.�H��۠jժX�x���͕7o�ѥ�/n	?��:��"iC����E����mWW���^*�cݺ��v�ߨQ�V�苺u�.+O.'2~66�@�PB.W���5k�E�FQ�^yԫWU���X,�f���F�.kР��mcc��%�`�Ӑ˗�o��4��}�����۵kO0u�/��c0u�+F�l##���P.W`�0O�>}2��^L	d2
%�͍ak[ӧwD׮�Z�6�n�x���7���`�:���'"""��I������i3i���Ɣ)_]N����Y���{�u��+��'�a��6z���IK6m�J�Jd�㕚*�B�v�#)I���h�8�6�̳�}��Ē%��.�����t {��,))ݺ��\�@P��`a��J=z3f�CJ���wG�ލ�.Im^���W_�����P(������/�֋�M�ￎ��1~7��Z�r����H@�]S��J%<<v���w8xP�^TTf�ޏC�n�W�F�?��^��([�(��G�[�� D T���D�9���<��=�ի��??%JX�gφB�DDDDDa�S�u����[���B��kJ�>>���OA(Z��v�E��Յ.Kc4p��51q�7T�cK$bT�T
C�~���
`��6������.�.m�-�.�������X�c��bŊ#�?��^\?z�
�z��3�b���8yr�A�t={6Ą	�TNT�P(����o������.�f��.]�c���q���� xM�<|�.]~A�N������.'W�R9~��8֬9GG[�\�NN�.K��J%���ɓ�f̸id$A�n��ڵ>���������5F�j�7KH�r��{���MFŊ%�.�������!����ѡ��(Y���MЋ p�z�M�œ'����=Zg�,���Tt����T*���	.\��ҥ���,ņ'�~�q�/_�D˖Մ.9W��Rѧ���$ (h��\[HDDDDW8���D.W`�X/�������Q�ǧ`֬���m-J���ɓ?`��v�6����	||�d���Q��5 ���S�|�ӧ��r�R��o#F��ϟ���\377���H �Сې��*pEDDDD�-��+����c�9���-����ǎ����{��,����ЧOc�K�)!!���3�dzO���ٳ��ի8L��q���|��F�.kдiel�:���y�t�pF���V�G�~M�.'K�^��ܹ�q��M���t�н�J�ذ�֮���6X��ڶ�!tY�:>n1m0sfg��!""""c�ˇG�^�S���޽�.�#t9*)�J��}?�3,]�G�È>y��-��ġC�СC]��c����,�/��xq/�[������!/��&갲2���D�����kL��W�>��{KL��Q�f�g���������[L���Ƶ�����e��~�q,[v������u�.�����4�!/�Ǝ����8z�;�)ST�r>�>��_��jմet�ZAC �ʱu�i�^}�JYc���pq�-tY*͘���W8	u��""""� ��<ز�4~�� v��s�߸�S���z�2���pq�����uR�nn����k<8Y�NTQ�1����ˏѧϯ�>�Əo't9R�t�a��q͛;b��>:,
���C1k�>�����qm1qb{����=� ��'���L������H��r!*����g4n\[�ՙi���3�"11��uC߾�u���N&S`۶3X��O-j���
]V��/cѹ�T�R
��ct��R""""���H�r���+bbp萇N�z�~�s�����`��� �@ɒ\AEE�᧟���ڴ��E�z�LO�{/ѣ�Z��:a��B�CDDDDj"�?�|���e������g�8�-+��KJ�{�\��a�x�66Ʒ�~ř3u���):vt_VŁ�X��/��HѠAE�{�J��F�jvX��0LL�ФIeA�!""""�`O^6���c��i�Pt�Z_�Z�<y�i�|q����"����TК(od2~��V����f�7�:w�'tY��:��3�aÆ����Y�r����������k���B�ލ�hQ/��J�ش�$V�>�J�J����~�
��C���{,^?�kh��������5͛�?��?��h��A�Z�����`�THN��K�5�H�
�,ذ���p|��<y�_cܸv\��\��3g�����5�5<<��wV.W`�pOܾ����K+�1�<�N�EP�M=�*T(���R�l�al�~͛W���}5:YGDD.]������D��]����H+���
��yK����	���&ؐ���$1'�ܜ�z�#��O��w�&���s� S�?~3f�!>>Ek�"���cǎmC�����{��Zm3&&�Ğ=�ѬY,^�ժ�i� x��:w��W���p.�AD�����|����"""QQqHI�!11))R$'K���
�TSS#��C,���ffF(Y���6(Y�
��EP�lQH$	C�S*�x��-BC_!44
qq�HJJE\\R �+acccc#XY�������Q�B	T�\J�I�H0�e��a\]Wa���7��Vێ���ܹ���nݜ��=P���V�vss x{{k�=]&���퍁
����O1k�>���s��
S�|kk�.�q�����+ƌi��3;k�m"*|��q�z������0<|���w��  #���������011���1��M`jj����'�+���)^�~�����6LM���h�j��P�F4iR	��<`&�S(��u+ǎ��������H$&� �����&��1���	$1޿OFj���)��|�7o� ffƨW�<5��֭��/���e�!�T���������Vk�J���W�`A ,-M�dIo�o_K+m�c����!H�B����e���X�ٳ��gφZ�U��ɓ}�~� ���Pk�Q�p��3��_�������+(�@ժ�ѰaET�Z���P�\q�����M�ڐJ刎~���8<y���G~��O�����	7���-��[7g�+WL͏�
���l�|
AA7���{T�Z_}U5k�E�j��Z�VV��?111�w��]Õ+�q���*e�.]�1|xT�\JÏ��C��p��]=���>��¢1m�/.\��{K��CGA&�`���.��t11	X��0��/�q�JX��j�,���/>�͛Oa��oѰaE��KD�)*����n�ѣWpt�EǎNhҤ26��Z������q�|(�����x4mZ}�6AϞ��G���������2e�bذpu����""b�ݻ/���7�ڵ>�M���%A��!��=W0e�n���(|�UM��'�)�i�I�Z�*U*��+���Y�e���K!/]HHf�ڇ[�"0thL��66�oW�P��};�_���(_����$"�������o��G�"�ٳz�l�ڵ�	]����N�������С[(Q�
�&�`���{�'>>�0o^ ʖ-��ۣ{��]�P"(�&V�>�g�b0gNWҜ��Cރ�pu]�#Zj���[�"��w����k��_cܸ���0��GC��!�g�e,Zt�3gv�ʤ<II���y %��'i�L;�7�B�M�N�_�����&�����ab��ً�#2�֭;o�pp(��k�P�^y��"'��1i�7��nb��v�:�U��vR�k��ڵ�е�3~�e ��*�
u�KN��S�հ�L�O�o����Xq��gѴie,_�Wg�O�D"T����6��Ő�...	K��ΝQ�~,Y�u�h�l�˗�pu]�z�*`�vw^�MD9��M��ѿ�ʕ'�<��G�l��x��-��n7.^���0~|;�K"%�+0q�7N��O��h֬���\��Æy��/�b˖a��.�
�_~�� <�k4��8q��-Ǟ=W�bE_���י��m��<)���~'T��66�X��7���H�~�̙{��]���,S�(�o��g`ɒCk��Û7���m-�={�#G<���^< ��/�ݻ�b޼nX��0.�$�Q?�t 'N��?�-x��fͪ`߾	�t�1V��K�rH@�6�9r��~+W����f&Z���Ǆ	;1h�8;;�̙��߿)�IS�թS���j� >�/�\�KP(4�4p���}�a�	����HD����R1`�&Kp��d�N�n"�#F����C�u�i�_\�H�\��۶��ƍC�[�S�k������v�߸~����@
e�{��-�Lٍ!C��s�zj����[/��ˏ��5�6�ںw�"�2��޸��3�&�޼�o~����e՞��D�۷1Μ���=b�t?t��nEh��޽a��6���=k���ۂ���I��=�P�����E�u�q��Xq!!��4r�����3ڶ�!t9�i۶�����*t!O.W`H     IDAT�����Ȃ�aa����Lم=�ԩ�pq���v��Ʋn�����ס�Y�/�m��2s��c����011B�N�1m��G�ˬY]дie��oGtt���OD����p��y˗�E��8}�>��'tYjѱ���m�3�
]
�3g��^`ƌN�J�p!G�������.�v-�χ
]
	�`C����0o^ ޾��@w��?q��sl�4��&jkO&S`Æh�n9���#0p2.��.��:BTz@��r�����j�,�}�&`�Z7;v-[.��_P�N�D�M�����#Fl�T*W۾�H�m�xu����ah�p؄���]����.�}��\y,t)�v�{�b�5k�W��޽ňۅ.�#��EФI%8,t)$ �y��W�u�i�j�g�>  �?���c޼n�^�NmmݺW�UX��&Ov��~��Զ}���Ju�O�m�3�H��=��ٙ�ׯ1f��W�Uj�occ��~���_�6!!!{�\����p��s�_��� ��.S(W�Z���]�.]
	 >>�uӧ��Q�8x�^�x�'�!9Y
 :��l�v�p�a��S���b5�P(q��} �۷	��F�l�#Gn�յ.�i��������}q�Ū�Cbb�eΠq�J8~|Z��5�S��A�j���1襱�2�ܹ�пS̚�]��A�~M0kVg�(Q��d�U�úu�0|�'j�.���[��j"�'.��?.����dr " ʏz���է	u���Tʽ�7�ѱ�j ���$�5.�|lR����k�I�ʥ��y,RSe:�F%��A��ݼ�w� �>�R�;�B$�`̘�������Ь�B̝�r��S��]��ص�2�.탽{'ڀ�S�Rw��jx��V�~~�q�`�>}_~�;v��L�(�]\jc�TW̟�8ޟ�0��I@�޿" �RSeP(�P(>�\Q*�Y�K*W.���h�� -333 �Ţl/S(VL�B��](�J�~�^�RH�2�>}�ƒ�~'�)��e,z�\����f����a&ON[�����y���͛x|��8p3���q��ج���k�T]G�y���y}���_vu��vuƙ3�1xps̟��W���'��I�ѡC]�ㅈ�5TJD��xqK��b�AFd)))���2|5j��o����w�X���2ꖒbX��{���矷U�i���J�;�]��ūW��Ո�KƐ![!���}�Ę<�r�~~WѪ�R\��^^#�e�0�.m8��U����mS ��ONm��M�� �!66/>��IH,-M1kVg?>ŋ[�{�u�<�QQq�ާH$�/������DRR�+&"]6gNW�iSFFYJ$&�g�۷	(^�R�2H _]��5����/��ur�fRRZ�+V������Bޛ7�����T*q�zΞ����'O�����/H���Gb�h/xx�B��p��a.�����2::׮=���U,_~���
T�6�j�B�^�q��-��̕�UKc��زe(.\E��K�u��|�477�o��īWq����U�BB"cÆ!�T�d�Aϐ\���W��=P��5$��_�"�E��^���(W�,,�7�<����̙����3��$�HDX��z�j�Ѷ���ر��u�+J�8��l���4U�^�tM:C9��H�q��+��'���A""b2�F��"�]t��c.]�F���S�zh׮&֮�a׮�X�����J��eo_7����y�i��F��α�1���(���B||
���O��
���&!!�.=ƪU��.�bii����G�u*�*Q����k�ɭ[�_���e� ��S�ǎ��r6L�D�5����i8��G�N���e�g9�Z.W��Ω�^!(�J<~���_ǜ9��}�H�����K}T�x��?�ڵ���ܿ��p#�B��T����ֵ�v�fnn�~�ӧ��l٢���WL��3_C8[�p���]�hQΝ{��j�HU�X;v� �z�GB�a���++S|�M�K!5n\	&|�ى�\�B^J�'O����k	]
	��B�B�����>v&�!�0aB;:���f������1�e����<�!���5*::ǎ�ŊG0p�fԪ5-Z,���.\�33���5�2+o���y�ҐHD�Hr���+W��f�L�*V,�?�����q�ZZ�X�M�N��:�1cڠS�z7n'�?��j�H�4kV+V���IHH��M�0bD��������pt,�QГ�:7\�n#%E�Qh��A���7���}�G�36��T)+��;ӧw�lV��d)�ۆ�Di�z�&M���铓�Rq��cl�|
c����M������`�(a��S;������å8|����!No\A(I���G�|gg�D9_�v��%������}K�}�M�>=cƴ�������=��>V��ҥm0bĎ�b�������G����#�w}��O ��1lX�K!`l,�ƍC?9�K=yJ�k���N����$4�A]�w��?�T���СC]�X�66��x?�������tB"C$B�m����$��/L��x�0
7o�#887n<���/!�)P����пS8;W��s�;ä���)����Ɯ9���MTy�	��z��KƔ)�!��aii�:uʡn]{89����=�T)�7פ�����;�w�F�7/ }�n@׮�1wn7�-[4�������s8\]Wcƌ�X�z��&"]0{v<x��gf���Yw�wf�S���Ν�m�p���`��T�n�Y����3N���욇�����شi�Х�@*�=zR�FF��H�dIo���8��{y����5 ����H �)�P(akk�/�tD�&�ѤI%T�f�됧P(�k�%L��ѣ[c���yxx�"��O��7��������n]{�hሉ����ʗ/^��(��{�pq��_~9�M�N�\U*�����I�J��ߗ	�����p�Z~��RSe��0A���2B_ݺ�pt����W�bIxy������s�Ѻ�RL��1c��NTŊ%�a�`�NN�>����&"!I$bl�8�;�Fh�+��)�{�^b�X/�����u�.�t̨Q�p�H._~@wz���S0o^ z�jGG[��!���2k����Q��\ @���q�88�����O�ǀ�  ��O,�r�Rhٲ:7��fͪ��.��ܹ���w�<�B�Dժ�q�̌\�?..!!�q#��Oq�f8��� ����h����z�4p@��e
�K��� �����>�H$���7�ٶ��hL���a��_�D�wo��3�Ri��oG $�BB"��?/��"��yz����st��ɩ�SRdظ�֮����=Ѻu����/G�z�Q���G�&��P)邰�h4o� p���Ϯ������曟Q�J)x{��"�ҋ�h�h ��å��4�"`�̽8p�&N������v|�\���M�
UO�ۡd��HH����� �_�x��05���ԗHM�@j�����R��c[&&&HIQ}���$,[v^^� �2��I���2�_R�����C]ZOݣG��P(Q�lQ8;;|r逺u�ae��www�رC���g�����=�^�c��b��}��|�\[[/���e2<�DHHDF��ݻ/��,���	j�*��/�����.��O��g��66�!�X#:zW��S�hG���!)��աK��<�u��y?k�,,\�P�2�e���X�h��e�̬
�남��P(��.'D��n����:60d�/_F�&M�.#_LMM����^--����DFn�h;�ell���ɏ5���t����φk��� �͛����H*���h���+�X\@�\�q��q�;��R
J���_���x�.������L&ǝ;���\aa��zy��3���`cc'�
pu�ggԯ_���_{m��puu�x;�@"��s�����ť6Z����ObٲèZ�t��02�V���U�,��O����x�0�Co_Z����W���
SS��?'��[�ժ���r�����7O5�$9Y3�jݧ>���A@@��e䛦^����'O�]F�=y����! h.tT }��Ehh�ކ���Tt��]��k��6t��tGVߗY^�צMM֣��r�g!���HL�懫W���S"��v#**o�&��X�Z���ٹng�
�R�t�'uQ���ˣ|��ZoW���a�d��Z���Q�fYԬY���}��d
��Fe����g�����Ĵ�W�V�L���G��Y�>}��F��T*��/�t���0��U�[��E��������`P�h[BB
V�>�͛O}�F�t�̔J%<<���sԩcSS>��N�3i�Q�FԨQ}��M $�+�*c�gH�3��w		)'҇y:9��\n��Q0e����!�5k��㳜Z?3�\���T��JՑ��HĨ^�ի�e�+�+��ѫ�����ӂ�D"��i%��&""""mb�ˇb�:c�ȼOT���[��%e�fQ~H$bT�f�j��ЫW# i�w<~��6�����?�9���ծ���Eժ�ѰaE�*e����$1LL�T^[�T*q�f�6K�BJ,�j��hР���!""""-�鞼�m���ɓB����Џּ�J�x��-""b���1���ǯ���Č�>x�V�r^_�H�d^7�[n��|MhVa{~�{�yy.
��F���凶^7:�􅱱+�DŊ%UnON�"<��?�EÆZ��H�2X�K/k����_3gvƷ�~%tIy�ۿ�6_R��N��={�����>=���kO0Ԑ.JJJ�ѣw�c�9\����/�����ei߇����X�����v�%tI���k�!O�̌3��"�����7�?��x��u�2��QW��
%.]z�FBB2��+�>}c�!�HW��dٿ�:���RSeH?���K2�Gً��GP�M��]ŭ[�H�.e��ߗWV8�%���<��m����t�en��e�f~���>D�ݧg��9����_������~���i��-;�^�GPP0���"$���%��� �����077QK[���s����s���
�֭��޽���M<���{ns3ӱ.����5��~y}�s�O~�gYm����Ru����k;y�ɩNu=�����~9m�/�B�˗# ���o >>FF���>���`���矷�w�5\��"�
�J�2YZ�JY��-m���9��SA��'�Ӏ�98�g[搦�����G՗����~�dw��n��m�"..�߂��5\��b�(c�B�T�|����	�~M�գG�p��WccI�sj�������~�y�U� QUOA�g�U�˩��\ym� ��zN�S���o�~��ػ�:���t�Őދ|�MJ�Ǐ��}�����~8��[?Zi�������B^n{��r��������"C��eVg�5�e�]m��V��憙�#�u[���p(i=I
��×[���� (�Zkɫ[�b [h�z(@h�Z�Z���WL���\y���T�ԕ[���Hi���׹���B�:��.Y 妽�g�� �9���T��E"�������=��I����ŋ�3�����~�߇�cll��=�#$$IIRH$"�d�#*�n;..I'����@n�6B����5yم'm+�7"ݑ��O�4yИ_J%P�X'\��$��=�!N��7�m���qi�KP)>�ϟ[ H[�1/����PU�W�����	]�F�+0�j{�"��ʂ>off�q�ڛ���22aƌ�j[,-�]�F	��(Z��.=��9}8fN�={�1c�4UV��D�޿��YyY���J����H��qRSCM
�O������_�޽�p��}��.�W/+4Ò%��ݶ:������AkȊ��_|���Ş=W�QBv~�}ڷ���*����&h�� To�&����>+�\%%��E���TZ~~W����\�/^��j����Z�&	�^x��Ǐ�����q�pRRd.U����V��8|�CKU����쮛��,��U��Vo����O�f�㚪�r�A���g�!=�Rt�� �1�o��e�z�Q#�D"H$Z��5XffrL��Μ���'����P�lQ Ș���}�7���nC���J[[sL�披W���!�e�0��ދ�����/}}=k�nڵ�����a���h׮��$��3vB��4ғ��n�{�2oSu;u���OD�*$��mX��~�ݖ�6�hQ��}7�/��������{�^��̷�*艂�������q��S�������m�A=��_��<�����z_��Βg�y��6T�SS������q8;W��s̛�/>���7p�@0��R �Hb�����]�:�kWg�{��ÇC��wW�<���+L🾆�zj	y��Ff7\��Е��i�}"�\Ng�s~'E�Mݦ��rbgWcƴ��1m���k������2�		)iWӲ�[g�M��qÆh����wÅ�ط���������4?����ןz��֖�����#�s��m!��Ѣ�#Z�p�ҥ�p��=��G��Fj�a��~W�އ�U��h��!*�H[+�Ν� �'O�5ֶ&���(����*t��kk]<�B��/c�������С[ظq�W��D�I�ʥ��w���AHH��-�.K�I$b�lY-[V���}q��=�;� M�T�4�B���:�E�u����#Gn#$$U����N�=��E0jTk��aa�F�rń.�PЋ��ݐʼ��r�����?�7a�ѣ�x�4QQq���"���*��ˏ��uC�T�ɩ<���]��111��k]��������9mצ��t�9���)z�n�޽	]�N*̯��Kb�d��(4�"䩻筠�+R�ʖ�oV��'�B�T9]�Pf]�_�wD���啦����j�N]����>$â!Oפ�����S��i!N�����%�U��&K#«W�q��3��D�رG �s�0""""���|HJ��/�a������D�,�5A �V�r02�t��>QQq	���҂]dd��%P����$""""��OE�Z`��0��N݃�}	�"�.xcc#��ģ[���v��sT� �"��?���e����!*�D"J���#G����=������>>>��OØq�����r�!����+������u�Bj�L�uyr�..� �)p�B(�o?�L�%���\��������P^��51��[���؏z�BB"���{�D"T�XNN�5�ՇI<�acc��:����H�dy��`�m�Q`r���6����H��E����HM5���{�|=]�S�N}�;�X���[�s��X� ��72~L�P(1rdkT�X�C�Rܾ����~
_߫X��O @�J�2�_��Ա�����xPPv�ܩ�vt�D"��իag��̧
�>>�0m�/�7w�޽������s�o�����{��遮<Ǝm''{ԩc�<�ѷo�יN*#!�E��n���	LL�`P������P��C]���0p�@��(H�R�� *���� t���#��K��i~"##����\��|���o����NN�aa�}p�v��� ���E���H�TX[���<��V�Z�/�r��K�0u�����z��f�I��}�&���y3-��#66�Ä-e?���޾*UJC,V�Q���|||ЧO��W������;ۃ��ןb���x� 

��]��v�?�Q������X�ʕK�n]��)���)k�����~V*��H+��Y��Lg�W9�G*���R(]:	q�A��y��t��~����ҥ��e�Ka>iF�%�'Au�̙3*t���C���g!O_���P��T iC�,�!C�g�ɻw�h�l!޽K��%
��@Ӧ�ѼyU4n\	u���y��L�-[Na��?��,��sy:4%Ϗ�ɓ׸y3"#�ݹ�))2�ؘ�ɩ4H�Y�~����y����� ����}$��yQQqX�8{�^�l�����P����}FD�|6)JLL�b�T)+뿱    IDAT�1Բnݴ:++S�=���v�	f�܇��#1jTkxx|K����8p3�¢q��/n��j����
7�	y 0x��:ur�"�m����5Q����w��S�_ ��?[�D,C,Nk��Fpv���ͫ�Y����K�l���ŋX̝�V��cȐ�~�R�����C�_Z�{��
%ʖ-�q]������s<ό!��'����y+WAj�\嵖�1���Dx��� ��޾M�D"���3B]�����wҫW�xq����EG,\�������?���'�N.BDDD�-��c���C$��İ�1úu�Ѷm��ٻ�&O��qqJ�(m� <�?4h���"..!!�q#m��͛ሊ��D"F�j��_�!�ǯZ5�,{%��yg���̙��
���1LL�P�lQ��&"66�����sNN�Q�v9XX�h󡨅L��o���ʕ�����uC���r}�nbܸ߱f�@���H��ѧjv���kaƌ�?�d
��&aР-6������&�{7Bp�S�����&J��R�6��Z5;ԯ_Ac�!?ll�ТE5�hQ-�w/^�f�~�����ԭk�ь����z����[̚�G�ޅX,�2���ٛ:���M�37׿@��K�a֬��¸qm1i�K���{/��#F�d�#"""�A��@����ĨT�$6m��5�|�M*��G��	�P9$/�D"ƱcߣF�2Y�FW��
<x��7�f��=x	�L��%������+ppH��O�����1d��<	�پ2+U��n����#**?�t ��7ЦMu,Z�+c6�܊�KB��`gW{�����DC�QV.���c <=�B*�� ]"C,a��.9��G��EEš}��x�6Ie�D"�ĉ�1m��F�צ��Tܹ���C8N�����
6\S�u��zy�,�&&���ov����L�m��`ժ?Q��,�W׺yޏ\��С�p��K���wz��鳼M�����ʀ��J�r,X��]��ի��lmm�}��kyI$b��� ))II��*]�,,LФIe���6AÆo�����N$A�T~�/��Իw'��7�����[WG�r�>�v��HսRw�<�J��p�|(ڷ_���cԨ�8sfF� �Z�Ν{O��xDDDD2�k� �q�033Frr��*J\���g�W�F��[	tǜ9�� )J�%֯?�#Gncٲ>hݺ�Fi�L��8�g��)��Y�¢��I4�>�����x�0ϟ�f�|��5ڴQ=���z�2���pq���~�硙�:t��r?��O�Y%"""*l.䙘�e�j8q����32���H�E�z~�ҹ��či��d
�ѷo|�m{����g�ǀ�лw#̟ߝk�^�����9sO\�����mU�t����f[~�Q�bIT�Xm�|�M�P�ŋXDDĠn����T*�֭��z�Q�*e/��pq�]�}޻��&�`ذ�߿��*%"""��2�� >�~>�O"�fM;�814���+V�E�*�o�Σk<��_;�$�!�c�SSUEyM�j(jH� �JԐ��K[CHЪ!!DJ�P1+���=��h�/5�Rj��(Ni$;ٿ?���!�������eU���s_Ye�\�����$O�Bz� IחtΟ��õ{��մi�V���M�Gq�2�{-�������ߛL���5֭��u�\\L*[�WV��C�o�s�a5o>UｷY����#�१�����]�	���JI  �(���<���r7\�[������,�˫�-�"E<4kV�||��r�U��ڱc�k*2r��u��_~I����Hu��֒�(E���z$�O��W_]��]���'Kj���2��<=��fs��H99���f'M   ;�%���W�*�M���%J<���A��tӠAK���d������ȑ��ҝ7�x�1OM��Ykּ��g/) `����.����D������f� YYٚ9�S=�|�8����Z�0Le��Z���ƭ�޽'�hQ����h  �^8eɓ�f͞�$����T�^E͜�]W�\�ȑ+�6Nݺ�u�0��Z3��lT�v3��i����ݺ[���oi���t�~PM��h��m��l�;F) �z�ä��Qb�n͜��U�X�   xtN[�"#[hժA���z�1OIR��i֬�Z��;-_����rww�С��m�pyz��M�銊Z�����^E�ڳoyݯ�����K���Y�=�zu��1J��hե�����5�c��F�kW�j�  �u8m�+^�[V����M�("��ƌY��~:g�1�|��V������d�W
���;[u{s��s�άݺ�ʽvü��w�L^���X�.##Kӧo�/Lѱc�|�@͛������43WZ�E�훨fͪjذ��zo   X�Ӗ����ZU��ҀI�v�l�{�L&���H;v�R�j���u�"#���߯Xu{���ɻ-��뵼�c>�5g��Ԭ�T��}�a�^Ҷm�դ�SV��?3�(__o͜ٽ�Ζ  ػY���]�K�N]Є	�l2FɒE���G�i׮#z������XF�}�?��z���޽T��ߵk�hED4��.�#F���?����p��x�d   <�Y�$�'�4uj�-ڭ-[��l��^����G�]��<8Yݻ����6/��e�F����ԩ�( `�~��>��5���R�REm6fl�gZ��[�����$   0V�-y�T[]��א!):}�w��������JM�S�~W@�͛��i�[(��$���'��&M��`�N��V۶W�FO�ṱ[�+:z�&L�矯bӱ   ��
tɓ����*Q�G����mӱ�ի�mۆk�� M��^��3t� �-�ގ;���x�훨*i�������������?�����իW#���Ħc  �:
|���*���_�������㹻���7�o����֭�q�?W�\St�FLѹs���:H�gwWɒ>6��_/�g���S��&N�d��   `��IR��%�Ys�n�֭�{>��1SSi��NZ��+5k6U�wɗ��֯ߧ^����/���y�_�b��}}'ͅ��tWBB��g  `=���_�����]�+22%�6Fqq1�w�h��Qz�����e��I�ŋW�e|ا#G�*$$N|�ƍ+k׮�
k�oE�b���7��ر�JN��N�   ��� �$*�����E��'i���6ۊ�V�J�aڴ�����>����ձ�s�2��V�\�:�����4s��-JHة*UJiݺ��S�|��>}�6n�^����I  ��,l��G��S���ROQQ������<y�/���Vttg�����e�c�jҤI�2�=���U�^�|�b�h���4~�Zed�5rd���H..��ڵ�)"b�bb:�g�F�>>   %�rН?��i�!��昆[���K1����Օյ��С4���={��k��z�v*^�ې,�~{B��sԣGC��l.  ��������k��ڲe�ʕ�3$Cf�Y�fm����T�������V-cHX����>}�.ܥ���jҤ�U����IK��6mf�F%&��
   ��w��fΔ$�_�B��{|���>|���;�4th+yz���b�hժ��4i����5zt[u���������3SAA�����ի��
  ������ĉt�j��kkڴC���X��G_):z����h��5n\��Lx0�֘1��׿~V�5rd���43Wvv����w�qm���a��   ��d�\9?͘��K�hٲ����b�+��C;v�R�*�ԥK�-8�˗�Ԙ1�j�z������'Clx����cS�k�%%���  8	f��CL�F��o׺u��Q���q$I7~��cS��cф	վ}m�#��E˗�I�6H�ƌi�.]��d2ni��v��w�(11L-[V7:   ���w��sԣ�<;v^�7�����ĉ�t�5o^U�'wVٲ�Fǂ���Ok���������9��||���u�֭����#�hР�F�  �Q��ӅWԪ���\��/~ծvܳ稆_��g/i��6
kb�F�ŋW5e�&-^���֭�I�:�Z5�c�E�Q	!!�����F�  ��Q���ߟT�����k�4|xk���Ef�Y3g~����T����{���SN�E)){�Q��3&P/�\�n�f�:~�7�T�:�`A���
   X%����Ѱa+�hQ�Z��ft��:����W�Nj�� ��FK�[����EcƬ����ԧO��f+�Z�����ΐ���֬y]^^���   ��=��C�iӦ�y�*_�q���&'Ǣ��݊�ި%|4uj�5z��XN�+�<y��-�ZTRTT'=�ti�c�QVV��w��ѣ�aC�J�.ft$   �%�!\�fV�������"�vF$-�F��X۶��.]���w�T�ha�c9��3�L�$OO7��n{�o_��f�X,z��dm�v@�WVժ�YD  `���t���z��PU�gw7:N�֯ߧ��N��"M��QAA����=�ѣW������y�J��F������]���ոqe��   ���u�!�-���Z��[��o7:N�ki���jѢ�\�޽t��E�cٕ>ت2e��ܹ����o���!CR4SŊy��O����०�Ul�g�:5��  P@��7n��!U��paM��^uꔷ���ryx��e��j��I-_��>��3y{{�f�'�v�a~ٺu�F�X!���v�j޸f6�hѢ�
O�ٳ���{]4vl���������o��H�4p`��q   �OX�i�'k��ڼy�]�\׮�5c�V͙�}���N�R`��:x0M��}���,�L&�RS�~�����c3f����_տ���la�3w�~��:u��_��ٳ��"  P�P� ##K/���W3�vm�||<��t_Lӈ�����Lo��RnF��7�����)=���9�$WWU��7ըQVk�|��M�(*��*V���i�_�YxU��Vrr���	   ���g%iiպ�tժUN��a3s��cѢE�s���iӺ�a�JFǲ���l�Ёi2���r��Ť��+�oߦjݺ�A	Nz�
���Ž�re����
   �a�+)]��,�_Դi���s�\\L
k���G�R����C�\�/�it4���\���V������O�N����\���^��K����R�   
(6^��2e��t颚0a��z���T)et����c����9U�\B		;�h�n���:��p�bc?SB�N���}�b�Ο��֭���d/++[����'ҵre�ʔ�s  ����6��۫�t��_�g�)ct�v��U��N˗�_|F11�U��s��-[�+,l������u�U�n�z4v  ��Q�l ;;Gݺ�����O�:�v�w��W?iĈ:w�F�n�޽���1�5���Ϩu�d6g�9�'Inn.2�sT�����ϱ������j%%}�a�   �Dɳ���]�*]���-�;fddiƌ����B�>�wM����v��������ͧ���+7v�����"��$�9[..&U���֭�g���ڶ��%3(����~�)S6iΜ�
�et   �J�<��f�}�ښ:5��8����36l���?�A��+2��
r��22�T��I�7�quuUV�Y&�Ie���n��]���}���W/�cÒ�Խz��dM���z����q   `'(y6�u�~��'j��64���q����C���w�j��w-)R_��+d6_��l�ã���(I���I��i��:���_e�\�^ǌ���(#c>��[���W����[팎   ;�S1�e��0��ƎMU��%ժUu�#�)33S:tPhh�]�s�Z�<<��c�Gg6[��f���kݻw��?����ҷߞ����յk}����8   �3��|ЧOc9rV��re��{��ё����`�c�5k��;v^�{'�I��4y��2�w#   ���瓨�Njܸ���*-��q��N�����9*_�q�����+}  p;~J�'��.�=����V��t�r�ё�@Ξ��.]���������r��a   ��(y����SK��ӅW5h�beg���C(����Phh�
rSJ� ��x	   v����J�.����/�ر�Fǁ��|9Cݻ�SFF�RR��ϯ�ё   `�(yx�r��멏>�J�����c����f#����=�����(%e�J�.ft$   8 J�AZ���ѣ��w�h���F��ww*jw+o��^�v���V�>u��y-[6@���	   ��g�A��+4��\�o�=at؉����H���вeT�rI�#  ��P��IM�<�޽t��oF�y(&���lۭ�n�����N3tw���3ww��3,����Qd�R��yD��T���ё   �`(yswwU\\O�+���x���at��[��*h�^�-m�Zv�WGb�X4z��ڸ�{%%�U�:匎   Dɳ^^����W�Գ�|�=C����v�Y<[�k&N\��˿Q||o5n\��8   pP�<;��WDK��WZ�%��PYY�FG��;-�������ߩY���e��F�  ���ّ���ҥ���'5dH�S�Pݼ\��[�7o��Oߢ�S�վ}m��   ��Q��Lժ�������):z��qȃ�u���%��&&����k5n\{u����8   p�<;Ըqe}�A7}��犍���8y�-dw*e7_��.�т;5v�j��N�����8   pnF��u�TG�.]�ر�U�L1u�T��Hw�׌�ݮݩ���w����ؓ��whܸ�;6P   N��g���i���K2$E%J��压eY�5��o���k���տ�F�  ��a���=��k)<|������qns�%���܂7~|
   l��g�L&�>���4���й:p�ёn���'.�M��N��w�<   �%����j��WT�V9u�:W��5:М9�+*j�&L��  ��(y�P!7%&���'K�k׹:~�7�#�>��~�I�6(*���ß7:   �%ρxyRRҫ��/�Ν?��ӿ	�0k�6EGoԤI/�O�&F�  @@�s0>>�JN�b�
+8x�~���ёp3g~�)S6):��^y�F�  @a��[�CJO�C�:��d2iժ���W�*��=�<88�*�s+W�Thh�����v�3�jڴ͊�鬞=Y�   ��P��ٳ�ԩS���=�j�k���z�{���[�駟��α���S���V����[���[4eJ�z�hh�{   �����N��]:�R�RE��2@�=�it��b�h�䍚3�sM����FG  @D�sǏ���g�B��)9����
���ɱ護>�ҥ{������u��  ����$>�Ν?�SO��G�*oo�#fs��xc�6l�^��ժUu�#  � ��9�C��ԥK�ʕ{\K����K7m-3Ӭ����k�%&��I����  ����d~��BB�D	-[6@Ŋ6:�Ӻr���Y�~8�%K^Uݺ��   P�щ�
�P>>^Z�l��:�+���x�z���_~����z�2FG   $Q���ӿ+8x���]�bE�J��1:��8s�BC�u��5��P�J%��   ��bt ؆���V�$�Ţ�g���ߍ���9����rq1iݺH
   �%ω�,YT����˫�:u�Չ�FGrh{�W��U�lq�^=H�J5:   pJ��{��"�����z�c��:z��ёҧ�PHH��ի�e��hQ6�  �}�� ���Z�"B�����)V��ɡ���QX�Bu��,�#OOw�#   w��+ȕ+�ԫ�|:tVII�l�/)++[nn.2�L�]�X,z�͚1�S�RÆ�d@B   ��0�W�x{{hɒ~�W��BB�i�FG2��bQÆQ���?����k���������M��  �aP�
/�BJH�n��_�EJH�it$�$$�ԙ3%I#F���zZ�Eu��/��I))����   �s7n�8�C ���ԼyUyz�ku�t骞��\\n_�?M�  �IDAT謎=���D��\_�|��Y�-�+�9[!!qru5i��ըQ��   ��ᙼn��}z�խ[^s������ёl�l�Q۶�u��Y����}դB�\d2��Q�J���-OCs   ��\``-�];X?�|^m�|�����bc����37<I�('Ǣ�E=5~
   %�^�_�|2T���

��u���f��?����rc�������_�ĉkH   X%�$?�"Z�l��v���4fL�23�Fǲ��L�"">�NK�!;;GII_�O�/��   V�3y�����4l�rU��7����O��*���+>~���s����}7^%K��8   `]���6����y�P��9j��}�������Ys�~�g�sss���h��%U��G~�   ���<�յkf��v��,���wo���;�p�BF�z`W�f�i��={Q����^���23�U���Z�xF�[��/Te�   8,J�iӦ4|�
��Vllժ��ёȨQ+�d�����d2���Efs�J�*��mk�U�jj��I��1�   �GɃN�<�={����˗3�x�u��eu�X^M��Χt��С�����_���讀5W��U�L�����ꪠ� ����oP   �J(yPXX�������l�]׮�l�T���YI����t�s]�vL����3�W�V��!   `}LW@׮]Shh������b8�ɤ�W�   xh<�    N��    N��    N��    N��C�L�z   @�(y�W�7   ��(y    �D(yxh&����ܭ3t��n~�n�}���4�ݾ~��    G�a�x(&�I�����v��-�m�����ƺ���Y   ��Q���r�ۣ|�V֚}��  �����&X"	   ���`   0�����3u    �3yx(7?�w�3yw��f�J^�{��   gC��C˫���ڭ�?���   @A�rM<f�    ��Lʽ�d   0%�b   ��k   ���   ���   ���   ���   ���AZ�t�L&S��%I�6��   ��L��/�N�<�={��.���*((Hnn�.   �D�    '�rM    p"�<    p"�<    p"n��    `�Q&ݖ���    IEND�B`�