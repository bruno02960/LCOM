�PNG

   IHDR  �   �   sO�u   bKGD � � �����    IDATx���w\g�����jCV����
(DMbb4��D/z���KrILr��%9/���c((b�A�ې"E�u���X!P@�م����%[f�òS�3��DDDDDDDDt���������f""""""�j�`&""""""�f"�5�B��
��1����������vJK()�@q���()�@AA�C���i������qi�j���W�Ѡ�DQ�L2����U���, ��~��4�\n�\KKS�ؘ���VVf��6�����f��4���	���aee;;K��Y�����05�f������!�(�D�P(���-AvvrsK��[�;w���S����� +K�Z^^	T*�C�0������acc[[]�imm�\++3���`n.���	LLt�I$��� ��R��V��r�j-*7��J(j �Z�Ei�_�waa ��T	�B���
����_TT��r
���QQ�By�EE-��\^UDW��Ӗh���ZY�uk�li}��lm��Q]�`&�A��]���|df ##�HO�=���ǝ;%�M��`�V�tE_��6h��-[Z�eKk�ic{{K���
c;;X[��Ĥi�����w��U�\TT���2�W=��_���b��=|B����nm�6mlѲ�5ڶ����-ڵ�G�6�pr�G�V6M�3$"""��Â���T*���p�F6�_�BRRRS� #� ��P*uW^�rڵ����=�������ۣ}{{�kg�-�Ѣ��r�ȿ�q��/}�J��*}^^	n�.Dvv123p�NqUq-�Jк�+�i;�mkg��ر��[���2�j"jz�Z���P���j��� �����T�hD�VTT��
���}������1rsK����7����SU ���A��@*����..������prr���=��к�m��<��	����ܾ]���"ܺU���"df '����HK�CY���G����:�hgg��:�N~��&"CRQ�B||&RRr��Q�����VN��%�h��n35�H$h�J������Z�Z����=z�E��07�7�oD����2DF��ڵ�HL�Ƶk�����v����Y�>�K�V��������ɡ�ӓ1b�Lt�Z�Ebb��3����L�ť��@wPakk�6�֭�vm����U����jj��J������<dd --7o��=�̫�o-��бcKt��
;���Kkt��
�;�B�-�r������B�;w��)�t)qqP�4055�{ס�dn˖�01����R�vv�J��H �F�B��r%A��b��o��]+�7�QQ��L&��Kk�C�v����Ъ���5Q��9�EXX""���pvv@�nmгg[8;����)����2*�Z���>W -M�OOM����LTT�ж�||�1eJ_��߅8�Z,��Y*-U���L��e�-��q��-(j����W�vpumww'���ݻ;�uk�c�)**Gjj.��� %�RSs������;�}��nq''t��
..�н�#�us��Kk��&�'��_���h����SSxzv@߾ѿ�<=�Ѿ�=$��- �Z7o��ʕ[HH��ٳ���L�R���W<�l?L�ܗ�35���d�����]���-ƍ����0dH7XY��{�*����8w����Z`��ј9s��A�a�LM� �z�6"#S������܁V+������pwo77'��9�[7GEO��B��]!��|��w������,dg��v��x���]���z�;j"�ɕ+����33��z`��~6��h-Z
5""���Q��(��+1n\o���ܜD�D�-==��N���\����Ø1��P����[w۶�������9L�஗e��a�LMNY�QQ7��R����2XZ�V�Y�ӧ#�ܜx��]QQ��
��>񩩹P�4�ɤ�ܹz�j�^�t}]]ۣs�V<�CԌ����w��޽ЫW;���8L��np���J5BB�j�Q�Ĥ������dt��R�hd$v����F��X��9��h���*²e��o���o����`&㗗W�S�����$DF� !!j�NN�߿�z�3�z�3z�vb�AK��V5s�z�6�^��+Wn#99*�r�=z�E��pum��=ۢw��<�C��	���kñti��[����ॷ+mE9��o�9���<|��d̜9X�Xd�V�<���«���G��V�9����ގ�=�bӦ�����o2~,����~%#<�*�ï!..R���Я��8�߿ڶ�;*�S�4HL�µkYHH�ĵk�q��-���=ԭ��U׵�{wG6F��T���vF�w|�h�X�;�Ri���X���~ ��v�,@�ڼ�4>�d�����O�7nd��W�ť�n}���f�3<Ap��-�8q��W��I(/W�ť5F��#zb��n��5;*Q�yp���\�z��J��2���nnNpww��W��9\�M"��F�����'O^ǆ�0xpW�#=�S��c����0�+V�d�Wȩq]�tO?���׳x��!bǩ���?��1k�P|����qH$,�� ��ȑ=z�N]Cvv1Z��°a=0bD����l�Jt/�F�����#�����t����D�^���ۻ#��;�˫z�lgtW�����K`��Sس���ݻ��qDdd2^z�g���,%v2�'��.]Zc��Yb�yȱcW0g�:?�!�ti-vf2YY�8t(����D ���.1�'F��wwg������u��_ll:JJ��0��]YD����"�]���)S~ĺus��ӴF�
���ſ�Сwѳg[��ض�>�lN���`��͛���r�\���QH,�IT))wp�`��cq�R*���=�~~7�7lm-ĎH��h�����h]�	�R[[��
�>}:�];{�#5+S��kk3�����s���W���O�;Z�x���eX�z��Q� L��#��0g�P;v?�p���<�|��U9s&�?�.|GG[��P#c�L�.66���	�ŕ+���`�	���끑#{��%�T*2��B�Ĥ�ڵ,h4Z8:��ӳ���Tu[6S�#5I��9>|)��鈨�4H$�Q�,��>�,v�q�L"�O_����X|4ciiy���%@.�A�PC.�A��`������gĎXE�����������ޛ!�X�EFF>v���ݑHL�F��������%S1hPW��$�\.��Wxyu���C��i����4DE��֭g�l�A��2xx8��.0���wA�V�"�D�-&&;vD`������4h4Z ���	**T"'l8�w���ǎ]���ŎC�())�ׇ#,�2n�̅L&�D��
�;ykjj�֭k�"�IѧOGDF��`n�X0�ޔ�*�ݻ#q�L"��,1eJ_,_>���O���YZ�bР�4��yo�.ğ&!""'O^úu��h�pqi����`�@]ݵk����L��=�jm��5 U��?7�={��ի�ŎB�쭷�#22��qu�mA`ggx]�:th��׳ĎA"`�L�ڵ�ظ�v튄J���1�X�~ƌq�a��\۶v�<�&O���,)Q "".��ܹ�BY�-[Z�w��ә�?Q5.\H�Z�+*��U6�nJ��,QPP&vjdk����ߠ��5�
�h����j�d�gcc��R��1H,��Ah4Z���cÆS8}�::wn�>�ôi�aoo)v<"�kk3���G��;���I�*�W�>�%K�an.��=hPWЅ��� ̞=YYE���B��V_@PVִ�KJ�EO3��h��{l��=Z�`�ǎ��03�8;�fz"��
���Yl�p�5�~��U�Ջ��"j�LL��۷���W_	@�g-2RW@8���C!��ЧO'�C�tG�~�`j�]5O��˗3vj��W��Z�l HI�A@���1H��^�:�//A����m�M�sr���W�_<:�z),,���'�~�I(�j���@̝;�g���!..���Һ�!YYE8s&�N]Ǯ]���C07���.:�;��/����D��+_ƤI�ō��6�V*�o�m��^����b�C�($���Y�>}99�ն�0Ă966�jPLj^X0S���c͚�ز�4LLdx��x��t�����-�N틩S���Z�̙D�>}7��7�����!C�cذ��ݻ=[�P�faa��[_����Faa�CW�+*�"%kx��_B�.�ѳg[���Hlm-�b��x���վnggXǕ���HK�À]ĎB"�}��V��J���b˖3��5�k��¬YCamm&v4"jb��rp��u�>}g�$"7����<�+����{�[7��MM�ŋ��:�G���{�6jT/l۶@�`��T��������Y����D����~}�C�ڥ��Ǡ�\��(6l8����./�fz��RV�>�5k����o�13g��'��	��+Wn����8u�:Ν����r�oo�Q�t������bG%j0{�\������Q��={���a|��~��wg�~ss���)j��o���V��77�#)�[���E��bĈ��8��| v���J���ͧ�|y(T*-���G�ʊW����H$�����k;̟?�QQ7~G�^Ǝ�!� �ޝ�F�������dԞy��^��+ª�f�B-r�'��u�±|�� 033��U����}�s��zqϞ���g��f�W��!AA������-��yñh�88�����

�~��Wq��ܺU��-�1th���+ڴ�;&Q�	��9s��ر+P�5���;V��������ݻ=֯�'v20?�x˖�V+�[�6�H�H ��2%ƌ�#G�Ĳe�ĎC"a�LU��2����p��<�||��ڵ�;Q�]�|'N\ŉWp��(����#G�ĨQ�0p��A��#z��r%|}����Yprr@D�?ŎT/��JL��yy�|-[Z���F����?���xyuDp�a����}ر#Ǐ GG�R��b�L��+ſ���~�}�t��OE�~�Ď�����$v�`jj������n�@T_��J�9s�����HL̆��9F��q�zc��;p7�퍱��{��ŵk�Ď!��֯� ���q�*��P�S����-ag�|OX���S�N;F����c���P*�7Z{a��6�w]��ys��A����~������M���C���UM�K�͘V+`ӦS���`XX��Ϟ���}����f��/�������$����6�͍��JK�Ñ#�8|8g�ހF�E�>�0~|o��W�v���!oo�}���'�g�X��`�4G�(�&�H�Ŏ!���$ ��v�ܹ�?����C��� ��P�˩-A�C"Q�uIIIx�嗱e��.G_y�WW5�/9�W3��>���X�p4�xc\��K��`ƌغu��Q�D"�J����:th��s�c���(-U�ĉ�8r$�օc���СƍsÄ	n<�+LMk��4��MSX��n݊3f���޶mۆ�3g���*�!7n�9I�3s�Lh4�cԛ!��ꪦ�%�f��T���'�ׇ�o��8|�=��)~�"��dee��=1q�'�Z��i�Ghh<6n<	++3���ǻa�x7�h������#��HX�e��;QR��ҥ�aƌAM��5Q}I����}�t��!3� G�$ 44���N����??O������A��DDD�HX07��e��}���<�L?|���j�*���Ӿ�=f��Y����T��G/#88˖ħ��3&N􄯯�ww;.��&�ȑ|����6��	�ŎDDd4������ o�T�<y!!�X���.=�n�������r��w?a"""z�&�ޫ��>���r*��-Ŏe�m�n��YQÓ�e3�cƸ�o�!""!!�ؿ�23�1l؝:�O"��jS��Q�5���Q�o]>�������;E��X��ޗ@��ԩk3��8q�*6mz?�8��r-U�x�����#�J0p�>�l2Ν��A"��6��ۘ{��X�NDF&#44�Q�%���D�M�p�p.]�)v��X7EE�ض�

�Ď"��:V��&D��`ٲ�X��&M�²e�X(533�%H�k�nc߾Kع3� ���DNE��DE�ľ}�k��� �H@E�
���ؽ;G�^�Z�AQQ.%v�&�sq�z/���9���x�bG2:�g-+�2��̣��*յ[�NW�<k;݃��pմ���7�:������/aǎ�~=r�*�����4m�e4��~�����;]]?��ͧ!��f��w���j����2*=�oQ����>�qu�=����}�.���#���wߺح[�_^c����j-N���={"q�`**ԐJ%�h�01�B�6Γ��X�w��$X07�7�ƒ%�w�v8|�=t��J�HF�q;��V��^{���S���cS%"�����p'���J��;#p��M�d��/ U�Ʈ���ꦫ��^�v�!����b�!�3u���2�'�L�U_EQff�ￄ�?��Wo�W$s]l>��A@dd
��{/�����X��-[*5�X���wb�lĊ�+��{;p�`�|s<�zkLL�{�1d���w>����3kDd\�y �Ph�kW$v�ĩS׫�'���"�Q�e}_{���s�_5H6�~�.�_C}��]^C��/E``4v�ą)M�ս�.�^BB&�]�"��Ut�	c���(���<�v���`6R��iX�p3
5~��o:��ؑ��Dd,-����\�{p^�
�Z_�����ͻ�A�{_�}W�<�&��eg7nn�Tͯ�'���JE_���`j�^��&ֺ�VKp�dk;���Nf=�� ظ����#f���ѽ{�^�!�v����6��_�����bŊ�в��ر���8�HD��4����u}�j�v����UkG���@Ll��/i�f���Q�>�R���~61�A�R�j:SS���bBB.]�5����>H���U()�Ctߍ�]Q��s�V�۷��3>JX�~��f#R\\���چ��x���-��g�A}�a�#ѽ�T��?�1x�x��{;wF 55���~Ցɤ��c�FLZ�O>�U�i��4��MAc�����QZ���L��s�vE";��뢵�����mEض-����w�1sK�@���ظq3���={.���8�TZH$�ۋU�=�/�(9k����і%�q.f#q�z^ye��عst;R����[����������c�LԴ��@�K��x�����2�w��='����Ʀ�����tCl��t�5]�y����˨n���e>����tO�{����{����#""{�^�޽PT�0ꑏ��u��LMM���__��({w܉k t�sM�sSfǹ,��@PP4�~{;�ܜ�s�"8:ڊ�ɪ��U}G��r��|c~BD�Qۘ�l�����	��N��� �?��}�.b�ދ(.�뀽�L� �Km�����u���~�c��$�cC�$�g����K"�`� ��%K����kػ���B�����U����u����sO��Bnn�݁�*�l �F��RY�&���I�6��?6�߅C*0�F���
Ă�1}�@���:�ez�(Q}I���|3qq_a˖��4�S�XD͎\.Ø1���Ǘ���5V�zcƸh�#$S�li�9s�"(�-�?�)>��ݺ9 lm-DN�<�
��*,,Â[����g��'v$��G���
,F�7"jz�rƍ�q�z��泥��\�HI��|m5v��Z�!�b07�������������57��{���E��bѢ�HO�煴F� �����YkQZ���77'�#Q-�Iۓ.���.,,Laaa*v�z���А��b��m(�i���,ŎPo�y]l��bGh6�$���={'� s<�6�e""#�̏ۈ���,�d۶s�>}F��ݻ������L���되h#v"""�6�6 �_�5kN��'��w}8���G�^�O?��ܹ�ׯ3Z�0�����'���    IDAT�z,�EVR���E� <�*V�|�'�;R�P\\��2XZ��DdX�j-���Oa�|�F�ҵ<�+fΜ)v<"""��"���ǬYk��[�ݻ�o�NbG2jYYE�GppN��++��]@RR������Sx��[�@w��RE�����]A��L��_L����l��D�H�Pc��?�f�1������˗�xh����$no�-����m*��!IJJ�����1�HS�F�`Ʌ��;w�p���pr�Hw�������X��ҥT���1zt/��?/ 8x=6n<��]������ \�r����H�D�STT�͛Oc��(.��/��ѹs���kmm�s�w{coo/v�'�駟��O?;Q�U�1�m�����;B�������_J��>&�BC�p��+W�++3�#A����:��Wo���
&����#G���� ���ߤ�v5$�T��Rk,X�	%%
�T�ZN'At��li��D�';�?�|��r 0{�P̟?m��<��!oo�R)����vl���d����艵h�]�t;F�����(h�Z��4I...pp0΋g��������,�َ����;0m� |��4�d��q�j-ΝKDpp�Eff�������ϱ�ܾ]���7"::ͣw�R��`��E���H�RR�`ժcر�<��-0�H̞=66�bG#"""��Iv#��0��_8v-��+q�����"44��epum�^ __xx8��Ij��{��_}�u����*WG"�
�Z�� ���+�p�@4:th�%K���̌�H""��W�� ����ذ�$���̙3T�H)/����	�ŉW�T���S]���??t��R��J``�~{;�J�ꇛhK�XZ�B.7����1thw�d4ΜIĊa8~�
�ܜ�x�X��{��
Ua��g*�o���`Ŋ����%v$�������X�����?�`b"���=����jž�bJL�Ƽy둒rj�_M��R)p�?LGPP��+��z  �C�v�\.1=�ôZ��aŊ0\������b��q5�'[��CX0�QI���oĥK�ذ��M�H���L��С8�Ʀ���c�􆟟F�v��5A3$eeJ������[�L���~�f�z�͛�
�FPP4��n�����������=X<��T*�칀�+�"11&�a��q�׏��#""���`֓��b���Zܾ]��[<t���D������n����GG;������C�tc1e6n<��>�W�<;:z	Z��~�ഴ<F���hDE����������ƈ,���)�u�Y�Ys99Ř2�/-�=ڊ����� f=��,��ϯ�V+`���Ͳ�B��ɓ��Ç�p�N	�vm__��z�O���J����\�t�&� ss9�����4iiy8p AAQ�t�&lm-���o�ٓ�3�E~~)6l8�NA�P��a��Q��=�	�v�f.�~,-M�c��j���#,�2BBbq��e��*���~~�"�{wG�#RP*��k���|8���(\�x66���q���F��	SS�JLO&3� k��֭gajj�y�c޼�h��J�hDDDd�X07���<��J�li��~[�����U�C���3g �u���'|}�Ѷ���	�Ped����F���T�ؘc�7x�x�:�~=+WŞ=Ъ�,��3�ʊc"Q��`n ׯg���W���۶-����ؑ��ƍ��ȗ.݄��cƸ�������������ܺU���hF���XY�a�wxa��^�.����T�X�Ç�������3��cS"""j,����Vc���3����21}�*����/��
s�� ��JCpp����Yh��
&����#F�dAC�֭��}���++3��/���� ���+�p�L"���ŋ���ǝc#Q�b�\Kg�$��~ ����)�Ĥa���pwwƦM����T̘F���ܹ�AHHn�.Dǎ-���__���2�T���ݾ]x��s4""�aiiz�x���ѽ`n.;"5"�F���bE��20rdO,Z4Æu;5Q,�ki��U8s&��˗�@�έ0s�������3����2%���u�H������TU$7�[c����
��<�?�KKS����<f��ѯT3�R�;�cժc�y3�&ya����p;5q,�k�ʕ[;���룒@*�ti��]�`��9F�_.7���!$$��W�Vkѿ���rGǎ��Xd����p��VU��S��^;�7�gw�t"v�8�￟��[�W��_��矏���Ӧ��믏F�.�1-5g,�k�7�b��KP�4�=/�H��S0��F�t��M���uo~�f.BB����d��H1bDO��y`�x7�li���D���]|_�lff�q�z���cǺ�k!�	����W �/��i��?����b�[�͛OA�0k�P���8:r�}"""j\,�#3� ~	�F[�{>�$ ��>�Q�+��G�������N��j5]||F���		�����ر������1�M��55o99�����h�={���ų��3���:v�
��Y�FAХKk�<�$�@]���X���o�66�x��;wX��� 6̏��`��p�՚G���WG�/��5Kbb6��[���;�h����ޮ�����'�СX������\�mk__w��ybР�Fی��6��)���\Y<��
/���⹑���c޼�j��k�#��M����?����(�o�F���i=���#����3TT�j������T?��ٱ�<>�p'�Z-�j��n�D���/к� @�P#<�*��cq�p��Jѽ��������Pu%��9�ͭ,��q�L"�r�}}����Ďؤ���6A�p�.G*��S��HI��^��aѢ1x��>���LDDDԘX0?�O?��o����D
A0uj?��:wn���ʔ��]ص+��{�ZR���4��c�.��Bo�����]��i�LD�,/�����:LLd3�+���,�R``^���z�|�I ����<�GDDD�sT*�������&�ˠ�h1eJ_��\\�3b�+�0o�z��T�$\*��gOG$&fcȐn��󄏏�!����R���"00
�O��Q�z! ��ǳx~R��]��ſB�?�w/)����6n8"""�Z`�\������~����\.�Z����}��>z�z�}�9|�����`W��D�?������-Qs��_Y<G����J%��66�bG4*;wF��C���f$	BC�C���)Q�`�� 6l)RSs���U(x��|ѭ��
��R��w��w�2�#�/�H�j�,<����257���8t(��Q8u�:$����&��x~����������v��aú���_�k."""��b�\���X̛���tL��w��A�^������̟��7�����~~�X�f�^�5W��e	��'O^�D"�ȑ=��	�xˣ���|��NH$�j�,��2H$h4��Ƈh��.|֘Q����롂�ƍ�0a��o?���A�j�`n�+�d���cnhj�9��X�X"��Yt�������&�HϢ��1e�bH�QQa���[_z��̈́Ba��\χ��JU�J�01QB*��L��L��T��L��T�Dnn:���K̞͓DDDd8�ҟ����$���b�1��% J`m�СQ�������Jh�� ��  �Z��@�����*deA�֠�Bł�H����z~�!T*����Ďe0�J��%5ڷ��������\���-[��f�LDDD�ƛ���k���j),,_}���*v�f�o�;B����&v"""��H�@DDDDDDd�X0U�3Q5X0UC���ѣ����D��|�ر'���݆���B���(��o��_;�C"y�=��1-�N���"�Vkq��5��{Ġ�BAp��U��S�xDDDDDDF��
�{��Vw���{_=z�C�k�Gu�U>��|ꓳr�Ϋ���e��%"#S�o�E��s����%P��  SS�d�N$�{��p�s��깚�{���}��ik��r�Y��\vM�!"""2VR0WW �����.�T>�k��$9뛧������L��s�vE +�r�*� �R�Hl��� �X���q]�����.@�7""""c�(M����>���|j;߆�}�3/��˗�b��$%�<P$kj���T����zg%j�rs�HdO4�G��+0� }�*u]��"��������lhf��Z-Ц�\,[v��G��
	��ƍ����Y�������b��P��@dDDD��T���W��TMy�GYߤR /o^�[E��D)����cǺ⥗7BJ��)$$��GA���mS�G�-֗�\&�>QScP�շ�!ɪ�|����)7���/`ٲ�p����s��A�TC"�@��V;���%<=;4rZ��#.�
����4��˫�b�Q�m�e�35R0Wvu��{=n��ͣ6�M�����'σ�{0O]�YWr��ǻa�x7��)q�pv����W�;N���HL�k�}oa���ԏ+`k[�>j�u]fm�Q�������5��G�O:���]�S�<5�\�e֗��)�L�)S���������#""R�J���3�Hj*�{���j��Q�k�'Y&#""���`�dS���[bƌA�1cn�.������Oa��t;��ͣ�����G��������oum@��Ҷ�,�F�����Qͨ������R0�xm�E15o���LDDDDu#; �!b�LDDDDDDT�DDDDDDD�`�LDDDDDDT��ھ}{c�  YY2���ՀVh4� H�V�n	�VK����Ix�M��-Ai�׮e������x���1,[�Z���b-��dz_�F���Qm۶3f�;�}*�=<< ��p��a1���=T�01��T��D�����J�{� @"��VA� ss)����^�Ұ`&�377wXXt�O?��F�� s�P��W��j�@���iH$�z[��$	���+v"""��H�k�"#����� ���`ʔ�x�!�ׯS�/�ĉ�X�pJKP�5��F&�b�Wl�<�����hq�L"���q�`rsK���/x�ť�ޖv��o@@�7~��E�#"""jd,�ka��_�o�Eh��rT*�uk��s���g���ּ����U��7#""Z���4R��}7/�0��25wj�g�\�*���J�� o��{�K�ɕ�ë�n�s��Ƿ�Nc�LDDD$̵p�v!�
J���9��J���$�<�^~y�z�K�,O�����a��P h���+�J�-[Z7Ȳ��+�Z�ӧ�#00
!!���+���sU�ܹs�F��E�~��/�ҥ�A"�4ڲ�����/,�k�����=������D�Z��w�:?{{�'^��ӉX�`#��P�n�-�Hк�5�Z>>�������ajZ�XnDt�J�ӧuW���c��_
O��¤I�[$Wڿ�/��gŗ_Ne�LDDD$"̵T^����_#'�5}d�W�5-^ye��r�/7;�������x������������c�++S��
??�ӻA��5*��N�$:���Rxyu@@�7&M�B�N-E˶sg�y�7�����E�ADDDD:,��`�ދX����<��w��A���
X�<�}R��RD�?���  �u� !!q	��ٳ��H$:�;��<0a��$��Q�48y�����q(,,��wǪ��:th!vDl�v~���>}4I�8DDDD�u"&N����6�tͳ{�n��{��]�ٳ7�`�&�C�ҠW�v8z�j�[XX���:�c�.��B�>}:���~~�zٗ��T��_CP��H.**��w����$B�\i������x�	x�]_���],�����T,��Y����[������6Wnn	���-8u�:�����~���TT�~����G^^)z�hw��y�˫�IR��T��+���+зoGL��+���Ď���?��;�O?}�;݃s=,Z�+�����K*���D�%K���YC��|�V�ѣ�1p�ll��GY�����d���"$$iiyh����������A]!�������)�j�8qAA�8t�"��Jre�C#����]��K��K/;=�s=ܺU������6S2�C�v���ױd�̝;\Ą���C�b���L��Ybܸ���u��Ѯ��l�f�DA�T���+
����q(.V�_��������ڷ�;�#i4Z|��.��q˗���)}ŎDDDDD�`�\O�}w˗�n3%�H��31uj_�X�o�9�ٳ�`ɒg`b";j����V]y��L�\.���=��-�ĎH͘Bq�\Zz�ܮ�aɕT*�|s��c���s0~��ؑ�����,�멼\��]? ����c��U�E��7�a��.X�f�Q��)7���!$$��W�Vk1`@��z���;�w�j>
5�����h��ƣ�T����/L��i4Er%�B��^ۄ3g�q�+6��ؑ�����X0?���x1o�9��A�bb�0{�z�ښc����ܹ�H)�\i�G�^ơCq8r$EE�pss�;�z�n/vDjB**T8v�
�����2%�� oL�艶m���heeJ̝�11�����Я_'�#�c�`֣[�
0w����aÆy0�E�HOL�����D�"$$YY��ԩ%||t�����2��4C'�PQ��ѣ������)1`��0q����C<?�/��iiyؾ}!O2	�zVV�����+�I���>�^ v�#������X$&f�eKkL��__w��ff&b�$UQ�BXX�q�H<**T8���ޘ4�m�؈�A���cƌ�P(�ؾ}!�NDDDdDX07�V��e�bE^}u>���&y611�jаK�n��B�1c\���q�z���B�$��r%��.#((
G�$@�PW�'z6�"�ҵk�1}�j88Xa۶pt�;��F�w�E���o8��Wς���ؑ�&+�!!q��ٳ� ����������F��ꮬL���E�ȑ(�j��&�[�nݴ��J.�����յ6n|�'�������F��y�6��\�M�^A��bGһ��r��]FHH,����2%��;������֭������)q�H���v��H���ܪ����*44n�ȑ=�j�,vM """2R,�E��U���7����X��e��[�H�F�P#<�*BB��;wJеk�������Ј�dJKU}����Ri0dH7���$�lٴ��J;v�������i��Ӛd�"""���H�J5>�p'v��?�1��}�DM�F�EddJU����\8:����~~�2��r��1��V�ʕG��
x�q����D�#G���G/C��`Ȑ�UEr�VzLmxV�<����o�������c�,��>�/��O?���Y7�LHȬ*���2`kk��cu����
kk3�#6I�����߶ <�  1q,-Mk|I����
�±cW�Vk0t��H��k~E2�1��/���?���%S1o�p�#Q`�l N������s�X�~ڷ�;������C����I01�b�������	�M�lc��NÜ9됛[
�Z�D�իg! ����W�-��q��eh��=E��_�\I�T��#((?�8O?�G�HDDDD�@X0���̝���%X�f6��&v$���W���x�"<�*T*���\��S��bG4J�7�Ƨ�� �h�  �L__w�];��8|8���8q�
�ZÆuG@�7||ܛu�\�����N/�  �IDATm@||֭��aú������fRZ��;��������`��QbG28eeJ?~!!�M@aa\]����>>���p��<�J%�����V|���pv��3)/W��~Ǿ}P��oj*���=q��5����{T���M�Vhuu�f.^z�g�����/��W�vbG""""�Ƃ����U��a������w�Md��L�����D����СXdf����=0p�K�F(~뭷�|��FH,�cǎaԨQ ���̙�))�P�5վ_"��ݽ=��__�&}����t�&��Y��m�e˫pt�;�fu��5,\�m��a����ܹ�ؑ� ��IGppBB�p��m�ha������끑#{��\^�3g�ą�u��FN�O=��n݊3f���h���6(���e 01����?�<�����X,Z�+��U�f�ʊ��5U,�Xzz>^yeRSs��O/c�XW�#����"88�.���L�ѣ{��������i�̙3�I��[���7��vm8$Z��333AB�װ�`�{�_��?ߏ�^���z��X&"""j�X08�B�>��wG��w}��[�yo�:��*���q	�ũS�!�??w��x���h�����u���Tu�N"���gc�$/=%3.�_|��ן������ǈ�����f#�q�I|��~����olm-Ďd���+p��e�����(-U��Z�>}���oM�`n�����Y*�@*�B��`��>X�j����
-�G�^���7�[nQ�łوDD$c���055��5����A�HFM�T�ԩ����йsi���,�Y�_����| �����^\\QuK)@7
�J���<p��wwl���Ν̞����ش�<�T�#Q#2; �^��]����{XT����w�b��h��5��fW������QD���XkL��%�}$��T�j�`4Uo���(^�Vr�FCML��	�M�0��[}\2  pf���y���9�w�yx|��;�d�Դik�Ds�k���f�rY͚y������%fGi0v�����z�a>\���?/ҳϮ����23c�ov$   42�X�b~���Z��9M��_���?�>}�JJJ͎�F���'33W#G.Q�Nm��5��  �DQ�]���U�f�jݺ�:x�BC����f�\�aJI٭�Gc���ڵ�qj  �&���z������w7�С��e��#.�ڵ2=��-Y�O��o~.OO�D  4e�o�����~ڲ%Z���Rt�:%$����fv,�wcy��ˤ-�͇��:z~�q-����__����С<m��ƍ�ev$   8
����PR�H�\9I۶}��#�����c�=�Ţ�����GmJ��V.�u9j���|�H�a(++N={�	   N���FBC�k��8�4d�"m���ّ�Z}ݑ�&���ocÆ��L={i۶�o�ّ   �D(�n&0�_۷�(22X11����h�TTؕ����3�5}� �X�Z��6;   ���5k��^�wޙ����THH�����X�S�t�ƍ[���?VZ�D͚ʒw   8Davc<�}�f) ���D˗`i/��#G
5xp�
/i۶��ّ   ��(�n�m�Vڸ�y���ܹ��8q�.]�jv,�s��\7�~0Qy[]��;�j��5j��u�޽���-��H   pr�&�j�(:z�22bt��y�@99�̎�����z���U.�����Ps%%��6�]%&nU|��^=Y�Z57;   \ ��	���eg�Tpp�"#�����Pyy�ٱ�s��=�t��{�6lx^11��  @�Q���V��+--J��ѪU96l�N�<gv,��ef�j��E��m������A�#  ��P���q�z);{�||�iȐ����Β_����
���VM��F���ڼy�ڵ���X   pA�f�y:th����Z�l���ۡ}��+5u�ڷ���h@��;wES���_�]iiQ1��`  ��an�<<�����;�o�-р��g�c���sZ!!u��5��GY  ��0C��ӟh׮8��Kqq��_���Sp	6�]o��S��o�O������:u���X   pf������0����cǾR���}��X@����K
_�+�ӂc�l��Eo�c  �Mp3~�w�N��4{�EE�Tdd������޵�ׯ�ɓ'͎� ��6J۷���t�o�Z{��3�  �zg1�K#�J�v}��^�$�ժy�FkȐ�fG�w999ڱc��1��jUBB����̎Ro�]+���ڸ�&M�ٳG�ۛ��   P�(̸�˗�))i��������ܹ�զMK�c�	:r�P��kU\|]��ՠA�̎   7FaF�8pB/��IW��jΜ�=�gfGBa�ٵx�-]�O}�vQJJ�ڶmev,   �9
3j���T������9�ׯ���#�}��pΜ����:u�f�����n{^6   ��u��'���o�={Y/��������J�A�1C�W����w�k�vZ�t����͎  �&�:++�iѢ=Z�l���RR�Qǎ\�w�����7���|��Rll�<=�   �w���"��mԉg���;H>>^fǂ���Z����۩h��Ա�޽�ٱ   �DQ�Q/l6�V�������9s��~��B�)(�Fqqu�h�bb*&f���<̎  �&�zu�|�������Gԯ_͝;Z:�1;���f�[o��թӽJM����>�c   f4�C����+�u��y�i�JG�*!!]yy;Hӧ�\e   8
3˴Q����Sk�|�޽Tr�+0�+`  ��P���X��[ef�*1q�l�
��j�F���}�  ��(�h4�.ӎ�zR3f��u�f�B#���"%%m�G��gz*1q����2;   P%
3��f׺u)5u��_/ׯ~�o�:��7���Wo��S����c����p���ٱ   �ۢ0�%%�Z����|�Oj��[		������\��ke�˻p��#��W���Wj�^5o_~Z?c�5   \���x�-ڭu�>V`����kذGd�R��Qq�u�@EE�������v����\%'g�ܹ+�:���O�-�MH   ��N�����,ef����jƌ�(�ى\�xUc���Μ� �ͮ_���z��Q7�����cJI٣S��)<��^zi��115   Pwf8�ӧ�+5u��m�T;ޫ3B���dg�^��ѿWQ�e��WH�||�����|}}�o��?�����6���V���LN   �
3�R^���fk�֣�С�bc),�1yyy���),��Q����ū7˲$yxX��ǋ���|���nJH�C�gbZ   ��P���

���~�����������}5a����1;Z�p��y��{]�rM6���[��V�^A�93T�<r�		  ��Ca�K(*�No�uP6|,�Ţ	����}u�}~fGs[�}��""����L_c�Z�x�XED�k#�   �.�����}�C�\��������ה)O�[� ����Ç�5n�r���TQ�Ù�,��ti���_l�t   @�0�%��W(#�����'�*88H�&�\���9��<xRQQ+e�U�n�ٟ�M����';5p2   �qQ�����������������ĉ�5~����5;��ٽ�3M��Z�aԨ,[,���� edD7|@   �Q�Ѩ�_����4��������+t��5?~]��������U�㸫��Rm���$��C2�J��*y{[��c�]wy�eK�||��ڵ�ڵ��8�;wVxxx��   ���jӦM3f����pUT�b�"��J��^�v��>!O�Ie�X�d�|�ϯe�J�������%���    ��y� MKyy�$)//��$0����5~�x�c    5b5;      Έ�    �f     �0    � �ps���   �K�0    � �     (�p	�����o�~��U�ڪ�W���cT�����zoՍQ�q*���   p�f n�b��0�=�����'��}�#{uc�.kuǭ�X��omƩ�{���   ���a�˫ka��_U�1��ͬ�f���Q��u�6�9��q)�   h*�a�K���_w^6���   pf����Ev'���    g��l�3f�o,Q6���d���m�<���   p�0���z>����j����W�v'�    M�.��r�����W���1m���벭1~O   ��bI6     0��F��'W��#̼   ����FM�u   p/,�    �
3     P�    p��    �\�����7;L��;   \	�����O�ԱcG��    @�,��A#2C������fG�IZ�n���@�c    �Ea    �.�    �f     �0    �����f�     ���<�u���s�    IEND�B`�