<map id="buffer_destructor" name="buffer_destructor">
<area shape="rect" id="node2" href="$group__game.html#ga8aead8655bcc62fb760afdf2fe161ab0" title="Destroys the enemy hit by the pong and desactivates it. " alt="" coords="348,107,427,133"/>
<area shape="rect" id="node3" href="$group__game.html#gaff72f275b5af37960b3baee51f855041" title="Makes a game round, where updating action on screen. " alt="" coords="491,132,545,159"/>
<area shape="rect" id="node4" href="$group__game.html#ga671b58f5509a3a9fa692bacccfc32cc9" title="Receives drivers interruptions. " alt="" coords="609,81,696,108"/>
<area shape="rect" id="node9" href="$group__game.html#ga425ea598437d36368c0e136f2be75a61" title="Makes enemies down movement. " alt="" coords="172,5,300,32"/>
<area shape="rect" id="node10" href="$group__print.html#ga4316256507429b01e848fd72e5fdca73" title="print_number" alt="" coords="187,208,285,235"/>
<area shape="rect" id="node5" href="$group__game.html#ga02fd73d861ef2e4aabb38c0c9ff82947" title="Makes game initialization. " alt="" coords="744,113,783,140"/>
<area shape="rect" id="node6" href="$group__print.html#ga92978930f74831bae9a6d6f22d089615" title="print_menu_kbd_or_mouse" alt="" coords="831,113,1009,140"/>
<area shape="rect" id="node7" href="$group__print.html#gae91d4cbee2dab64187187499dd0eecd4" title="print_menu" alt="" coords="1057,113,1144,140"/>
<area shape="rect" id="node8" href="$group__spaceinvaders.html#ga3c04138a5bfe5d72780bb7e82a18e627" title="main" alt="" coords="1192,113,1243,140"/>
<area shape="rect" id="node11" href="$group__print.html#ga1243268c621c2049a41956ccfc934fd5" title="print_info" alt="" coords="350,208,425,235"/>
<area shape="rect" id="node12" href="$group__print.html#gabbb46faef7390f85ad76868944abcf20" title="print_score" alt="" coords="475,208,561,235"/>
</map>
