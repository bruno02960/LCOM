<map id="fire_pong" name="fire_pong">
<area shape="rect" id="node2" href="$group__xpm.html#gab41dd197773f68e69e18c73a8119ba5e" title="object_creator" alt="" coords="128,56,232,83"/>
<area shape="rect" id="node3" href="$group__video__gr.html#ga1cd7727ad0fc3fe3ffbbb98cd9115c1c" title="Returns a pointer to Buffer. " alt="" coords="283,5,356,32"/>
<area shape="rect" id="node4" href="$group__video__gr.html#gaa55320d571dc2cb8179422a9d8114de0" title="Returns horizontal resolution. " alt="" coords="407,56,479,83"/>
<area shape="rect" id="node5" href="$group__xpm.html#ga05b2c5e4dbcaffa701703b50a2111783" title="read_xpm" alt="" coords="280,107,359,133"/>
<area shape="rect" id="node6" href="$group__video__gr.html#ga36218c155eade74951ce7ffd60711a9e" title="Returns vertical resolution. " alt="" coords="407,107,479,133"/>
</map>
