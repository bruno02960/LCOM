�PNG

   IHDR  �   %   ���   bKGD � � �����  �IDATx���Mhg���n���C1hA?
Qhsp�L��J�!b�[�!�\$��G�x*�f7qC��w-i��lU�L��+m>4[m����M7���|�3����dg�}�gvw�gf�I�t:��8��3 "����BDD±��p,.DD$�O� �����d҉|H��M�p��q��0��'������ӧQVV�t*�9rcccN�!D��I�?-v��8p UUUv�F*��( ���e�OuuuN�BE$���󨯯w:C$I ��`�����ޕKF{{��)�V���8v��i�����t
TD2�����8fdN�p΅���cq!""�X\��H8""�(�Kuu��1��!33y�Ɖ_;r6Í�'����ϒ��!��H��%�)D"���=��'�N�qn}��jZ��`������itt\ř3�y�����/����tCC�����a��� �@`#����19Go�o�1::�4�>\�'��@Hq���F$y�VQ��}�:=g���)�/�7�6�r=��1���xf<x���(:;�����x�H,�%����;��3f�3����zI��m�y��\���:-�!o�+_��"���e�˼V�VO<��`F<>��Wk���,摉�q��b�)�g��{�֧(®\��|�����O=���Q��L�F�1>>�TP�>�sYA��t;��k��k��*�1��h<=mE�_���g������q������w�D
��Ri �D�0����3KXq�3`\�����|��mE�xJq�܏�q���^����*���K��������6Fs����mն��ӳ�"�!7	cco��r����ݻ9x�,,����@�N��i��̈��s��j1�[�g>fp���X��;=zyi��B���N���B[[�plQ��uB��ꉗ\����AS��+����}X��k�=�hٲLaQ35Ǻu-�㉶r���_O�tq��Y
�O���Z�JB<>�@`���WB2��{@J���� v��j8������ڧU��3{=�D����O��݇x��m���<��9�|���z�G8q�[����o�9��V���#��蜋��!> H0;�3��~���4zzFq�� �<y�ϫz�}�gػ�i6;{��;���>�����U[gt �b��f�5KD�D�/:�uu��>DW�0�]��D"	I��L*����1 ��-q������d�FoE����S�����u�Xѧ���k�ԴMM���q��(��ALLL/��w;�y3�T��]'*���y��*=y��W!�.,)񢦦55�x�vׯ�C(4��7-ͻ�R��h����t�����o+&�s��KD��b4�Q[����uZ[�`d���#������EQh�N>��կVF��KD�����vF�Yq�TZ�Gmmjk+03�W�,�����3x<�W3/_��z�O�IG�ߕ^�U�s.�_E�TTl@{�7�u�wtw����_\�L?�Y�|R����hh؉X�5zzFq��(/�p	��hqQ��U��^��y�TVnFe�f�:���t����7N�������X���*�S��8Z\X@�͊���~Paq��!"����BDD±��p,.DD$\�	�h4jc�K�|�`���
J0DII��i��v\Ki٣"�'E���~���9��!�>�Un߾�;v8��!+V������i�c|j~�����9""�Ņ���cq!""�X\��H���:gH�    IEND�B`�