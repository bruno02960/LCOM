<map id="round" name="round">
<area shape="rect" id="node2" href="$group__print.html#ga1243268c621c2049a41956ccfc934fd5" title="print_info" alt="" coords="117,107,191,133"/>
<area shape="rect" id="node4" href="$group__xpm.html#ga8b990eb150243edd20fb9c4182748528" title="buffer_destructor" alt="" coords="404,56,523,83"/>
<area shape="rect" id="node10" href="$group__video__gr.html#gabdd05df698103c4641478f491e11e284" title="Copies buffer to video_mem. " alt="" coords="393,208,533,235"/>
<area shape="rect" id="node12" href="$group__game.html#ga9a691a2142903ae9009a88a62464ddd9" title="Says if there are still enemies. " alt="" coords="108,259,200,285"/>
<area shape="rect" id="node13" href="$group__xpm.html#gab41dd197773f68e69e18c73a8119ba5e" title="object_creator" alt="" coords="411,157,515,184"/>
<area shape="rect" id="node14" href="$group__game.html#ga8aead8655bcc62fb760afdf2fe161ab0" title="Destroys the enemy hit by the pong and desactivates it. " alt="" coords="257,5,336,32"/>
<area shape="rect" id="node3" href="$group__print.html#ga4316256507429b01e848fd72e5fdca73" title="print_number" alt="" coords="248,107,345,133"/>
<area shape="rect" id="node7" href="$group__xpm.html#gac0e395e7e8c65b90f0680c7a917f1acc" title="title_creator" alt="" coords="418,107,509,133"/>
<area shape="rect" id="node5" href="$group__video__gr.html#ga1cd7727ad0fc3fe3ffbbb98cd9115c1c" title="Returns a pointer to Buffer. " alt="" coords="601,56,674,83"/>
<area shape="rect" id="node6" href="$group__video__gr.html#gaa55320d571dc2cb8179422a9d8114de0" title="Returns horizontal resolution. " alt="" coords="741,107,813,133"/>
<area shape="rect" id="node8" href="$group__xpm.html#ga05b2c5e4dbcaffa701703b50a2111783" title="read_xpm" alt="" coords="598,157,677,184"/>
<area shape="rect" id="node9" href="$group__video__gr.html#ga36218c155eade74951ce7ffd60711a9e" title="Returns vertical resolution. " alt="" coords="741,233,813,260"/>
<area shape="rect" id="node11" href="$group__video__gr.html#ga5c30cdd3eab0edd2734ab3871f7000c7" title="Returns number of bits per pixel. " alt="" coords="581,259,693,285"/>
</map>
