<map id="read_xpm" name="read_xpm">
<area shape="rect" id="node2" href="$group__xpm.html#gab41dd197773f68e69e18c73a8119ba5e" title="object_creator" alt="" coords="416,385,520,412"/>
<area shape="rect" id="node11" href="$group__xpm.html#gac0e395e7e8c65b90f0680c7a917f1acc" title="title_creator" alt="" coords="132,169,223,196"/>
<area shape="rect" id="node3" href="$group__game.html#ga02fd73d861ef2e4aabb38c0c9ff82947" title="Makes game initialization. " alt="" coords="940,195,979,221"/>
<area shape="rect" id="node7" href="$group__game.html#ga1fd9e64dab3abe9facfb4dd7e1267bae" title="Creates the pong and switches game state. " alt="" coords="595,347,669,373"/>
<area shape="rect" id="node8" href="$group__game.html#ga671b58f5509a3a9fa692bacccfc32cc9" title="Receives drivers interruptions. " alt="" coords="754,321,841,348"/>
<area shape="rect" id="node9" href="$group__game.html#gaff72f275b5af37960b3baee51f855041" title="Makes a game round, where updating action on screen. " alt="" coords="605,245,659,272"/>
<area shape="rect" id="node10" href="$group__game.html#ga425ea598437d36368c0e136f2be75a61" title="Makes enemies down movement. " alt="" coords="568,397,696,424"/>
<area shape="rect" id="node4" href="$group__print.html#ga92978930f74831bae9a6d6f22d089615" title="print_menu_kbd_or_mouse" alt="" coords="1068,117,1247,144"/>
<area shape="rect" id="node5" href="$group__print.html#gae91d4cbee2dab64187187499dd0eecd4" title="print_menu" alt="" coords="1295,43,1381,69"/>
<area shape="rect" id="node6" href="$group__spaceinvaders.html#ga3c04138a5bfe5d72780bb7e82a18e627" title="main" alt="" coords="1429,43,1480,69"/>
<area shape="rect" id="node12" href="$group__print.html#gabbb46faef7390f85ad76868944abcf20" title="print_score" alt="" coords="425,195,511,221"/>
<area shape="rect" id="node13" href="$group__print.html#ga5f04c1438b5689bedddc17eb0dd9d060" title="print_message" alt="" coords="744,144,851,171"/>
<area shape="rect" id="node14" href="$group__print.html#ga4316256507429b01e848fd72e5fdca73" title="print_number" alt="" coords="271,245,368,272"/>
<area shape="rect" id="node16" href="$group__print.html#ga2eb771fa3527f72e821a14e413498d1d" title="print_instructions" alt="" coords="899,43,1020,69"/>
<area shape="rect" id="node15" href="$group__print.html#ga1243268c621c2049a41956ccfc934fd5" title="print_info" alt="" coords="431,245,505,272"/>
</map>
