�PNG

   IHDR  =     $a   bKGD � � �����    IDATx���wx�e��ӽ�^t2�(�A�^dO��C�-***�@^e��P�! C���)-�Q
t�t&�Iw��B�W�>�s]�դM�I������6P��j�C��,=�������H'�� """""""�d,t ""}SYY��**jPS�DEE5�r%�j@*����S^^{""]c`` ;;���&&F��4 XZ������氲2*"i1�DDOH�V�����e(,,CQQ9d�J�dՐ�*!�VA*��LVUwY*�De�UUrTUՠ�Z!�� "�JFF���6������accGG+��������pv����M�e#�c���{�;�R�X���bde#7�����((�A"������P(T�}���ll,`kk^������氳����9��M`aa
33c���<v��������u�gl��g���ޞ�H�(�*��U�]�-�k⊊j�dU�ɪQVV��
���J�PVV���rH$R� K!��~?pw����4p���S�e__'�����c%"���҃�t�Z�FNN	���^���"�� +�����K��#���������pv����-�����dWW[89Y�����V044���#UUrH$҇�YY���(ăx�֭���4EP��4qG�F�7��8�����
�D�3��*��Jꎴ������ ��`//{xz:��������r���=����b�"��H��ť��(Dzz��Ÿ?���!+�j����h��M�z�U�	�Fp�'O�!"�R,=�H+=xP���$&f#))��9x� `ff�� W�  ������Y
����4QEEM]��,���ٸq#��055F�f�	�A�Vв�5rgIND�Xz����(D\\:�_��ȅTZ	ccC����Y3/4o�fͼ�//>%"��B$*�͛��q#		p�v6d�*��Y�MDF 22 !!>\BD��Xz�F����ƍL�ǋ��DKKS�h��`��%�7�4�7�""���R���*All�\�=23�`ii��P_DF�]���c	BD�Xz��*+k��s�����Tܺ��\	//DD�#<���~h����jBDD$���\��ZW�$'�aii��S�F��5~~�B�$"�K,=��^)*ܸ������ܹ���A�P�yso�k��� �n� ���J�����D"Ù3wq��=�9s��e��uB�΍ѵk0:th++3�c��D�ť8z4'O&�ҥH�UpAǎ�СCC�o���0JDD�G�R�Ν�:��3g����t�c�F�ի9z�l�c�,�D�Bܻ��#Gn�ȑ[HHȄ��9�uF�΍ѡCCxy9�����I�U8u*	���ɓI(/�F�־��n��_A@�����t
K"z.T*5�^MǑ#�p��m�D��v@���QQ��FDD�r�.$?|��6��JѨ�;h���[�ߟѳb�AD��Ν����{�!'�-Zx�g�ڢ�Y3/��i�Z���L��11	��-A˖>��?�����������K"zj��Eس���ǽ{yp���a4(��J=#�J���4��\���	()�@D�?E���9���)�� �'RYY����ض�
��Dpu�A�~�1p`(Z�j t<"""��P�p��}��\�o�݄\�Dtts����7�������4K"�[���a��ص�*���۷�G��add(t<"""�Q^^�n`��X\��OO{��C#���,t<""��҃��Ku���'`�拸z5���=�-�o�%�DDD@$*�ΝW�c�U�� 22 cƴC�>!055:��`�ADu$֯?�͛/�����-0fL;�k.�%""�4*�.$c˖K8t���,0rdF�noonOD�҃�p�~֬9�_����&L脑#���l-t4"""zBb�[�^�����/C��M��k�ѩSc�� "��҃H�]���5kN�ĉ$4l�ɓ;c��p.�%""�b
�
G��Ɔ�q�B
���1aB	kk3���+�DzF�V���;X��n��D��A�<�+�w�),DDD:&5U����c��+0661�0aBxx����^�� �#'N$aɒøq#���1sf�������^���
���%���9��_�֘<��7�:��҃H�9s_}uׯ?�K/5�ܹ�h��[�XDDDT��r%bb�c͚�HL�F��A�2��u:��҃H�]���ŋ���tt���s_F˖\�ADDD�����z�i�<���̚�={6��S"�),=�t�HT�O?݇C�n�S��x睗�+t,"""�@�ogc��8|�6tÌ=Я_+
��虱� �!EE�X��8֯?|�qt��D�XDDD�����ʕ's�ގ�>�;�������ш��5�D:@.WbݺsX��(�͍1kV/����|�������HT��;�;b��n�9sza��p>� "��҃H˝={���B^^)&O�iӺ���L�XDDD�岳��|�1l�~��Θ;7}����"�*,=���X,ł{s}��Ă���� t,"""�1"Q�.=�ݻ�Ѹ�;�~�e���,?�H�� �2*��7_ĢE�����}6=z4:��d1���0���ơ��;7:��b�A�E���;;p�v6����`Μ���0:�;wr�x�A;���]����_A�f^B�""��Xzi�����0֬9��P?|��4i�!t,"""�c/�������L��s�y�-i�D�ƍL̞�YYE���~=�-ϡ%"""��V�s��X,ŤI����`kk!t4"" ,=�4�\����G�r�qDEb��W���wO���H���J�[w�~{ 0w��=�-��%"��� �@w��`ƌ-�
��}��k�����4�TZ��ˏbݺsh��D�vAB�""=�҃H��Tj|��I|��!���a����s:�SIO�����q��]���O>�yD$�DB"�aƌ-�|9���&u��!Ww��:u�.>�p7rrJ0yrL��,-����D��默9s+��ͱj���������x4�c�򣰱1ǂ�ѧOK�c��`�A$ �\�ŋbժS4(�����б�������|>�|?v�C������A��u:�8�Dy�S�l���b|��`!t$"""���T�]��(Č/��7����H�XD��Xz	�ԩ��6�gxz�c͚qp:Q��˕X��4�-;
{,Z4:4:� �D�H�Vc����C2$_~9ff�B�""""DVV1��ߍ�GocȐp,X0 ��VB�""�҃���dU�9s+N����bܸ�BG""""�G���{����.��C��DD:��Q=HNc���(+��ڵ��/t$""""�"�U�/`Ӧ���=�����б�H˱� z���3��iS/�]�\]m��DDDD��._N��o�D"�{ｂ�c����@�XD��Xz�@�_|q �Ƶǂ8������	TW+�l�|��I���aٲ����w"zz,=�^ �\���ۅ��c�p� ��Q�HDDDDZ'11�goCjj>>����\�ADO���sVZZ�I�6"!!�W�C�n�BG""""�Z
�
�|s+VCx��-{8	���K��H$*�ر?��F�&�I�#�۷�1c�deᣏ�cԨ(�� ��҃�9��aܸ��~�ggk�#锚���0V�>�N�aɒpw�:i0�D���c�x�Mx饦��Q033:�κv-�fmE~~/�~�Z	��4K�g�m�e���N���jDDDD���J�O?݇.`��p|�� �ؘ��4K�g�b�1|��!���˘9���q�����ΉI�3g,-M�r�(�����4K�A�T���bӦ���aĈH�#魂�2���/8u*	3f���Y=all(t,"� ,=��RM�Ӧ��'��z�X���L�HDDDDzO�VcӦ�X�p�6��wߍ�ֶD�҃�iTV�`��q#�7OBX��Б�������Ř6�g�D�����ۗCN��K�'TVV��c@J���2M�z
��������>�d6l8�Q���駃����b�A�JK+0j�Zdg�`�Ω
r:��Çoa��_��i�5k^�s8"=��>D����C�~��|bb��K""""-�Ǐυ�����`��X�#Q=�J��!�bذUP��ؾ}
<=텎DDDDDOI�Pa��X��$Ǘ_����б���� �99%2�;�����_����F�HDDDD�Μ��i�~���֭�#���[�������������&""""йsc><VV���^��~�!t$"z��҃�OrsK0x�w��4ŎS��h%t$""""z��r%,����1iR'|�A_��	��^ �D��W���kOiٱc
�����DDDDD/HL�u̝�͛{aժ�pw�:=g,=��kSSc��9���HI�`u(-��ڵ�!22@�HD�q� �X�!C����""""=�C�� **Æ}�.���#�� �WXX�A�����v�z��,<�����Z��wߝ���1lX,Z4���B�"�g�҃��TZ�!C�EYY5��77[�#��N�Lo��� ���x�� �r<���VeeF�^���r��1���[�`:4ee�x�奈�K:=����r%^{m���k�Tx{;�����4���3���0?��o�:�K<���B�����˗S�g�t{�����4�Z�ƲeG�d�L���������б��)�� ��T�0s�V9r۷OAh��Б����H���\ǬY[ѭ[0V�KKS�#�b�Az��va��Xl�4	:4:i��xƏ_OOl�8nnpJ�8Ӄ���_��?_���cYx�S	����s �+л�r$&f��� K�7^��eG��W�гgs�����v@L�L{`���8z��Б���� ����ߍ���#"��CDDDDZ���7��a��`�����BG"������ΟOƨQk0n\{,\8P�8DDDD�C~��>�x/�k�E�����H�HD�',=Hgݾ��!C��K/5�ʕ���=wg������ ?�0vv�BG"�?`�A:I$*@߾+м�6m��֝����^�{��0n܏055�ƍ����E�HD�gz��),,�ȑk�����'�� """��qcw80vv���g9bcӄ�DD�� �RYY�q�~ l��:,,LNDDDDD�����v��N�cĈ��مHC�� ��T�0e�fddb���pr�:�33c�Z5cƴ�ĉ?a۶�BG"�{�B z^��ߍs��c�Ω��s:�!|�� �����w@"�a��B�"�[,=H'���9l�t+W�Bh���q����HϽ�fw8;���#?_���А�	�7�������>ڋ���A��CDDDD >�����PPP��+Gq�>Q=㖵�ծ]��С�cذ,Z4D�8DDDDD�%>^�1c~@���X�~��̈́�D�7Xz����-AϞK�u���Ȉsy����H3ݿ���#�����7O����Б��K�J5��w9  &f&�r""""�x99%9rjjض���:	�H��q�:J�
S�n�D"æM�Xx�V����޽���d���W 11[�HD:��i�/�<�S���q����r:����ĎSвe�-.\H:�Nc�AZe��X|��I,[�*��%""""�daa�u�&�w���ǎ%
�Hg�� �q�r*�yg�M�έi����H�b��?�^�'�ߟ t$"�d,t �'!`Ҥx饦�7���q���������>��?��M0u�f��(0xp�б�t
K�xRi&N\OO{|��h������y��ް�4ŬY�PU%ǨQm��D�3Xz�F�ݩeJJ*q��LXX�
�����蹛>�%����ww��F���;
�H'�� ��`A.]J�ΝS��a/t""""�f��.077������J9�N�&t$"��҃4֦M�~�9�Z5�;��^7�=��M0w�vTU�1gN/�#i5���ΟOƇ��[o�B�~���CDDDDTo�o33c̘���r|��+BG"�Z,=H�<ک�WZb��B�!""""�w����o����r|�� �'��j�Z�D�H�U��^GG+��9��K����H��8��I�~�СX�hY|=C�=�T�0e�FTW+�~�DDDDD���wƦM�c׮8̞�J�J�HDZ��i�ŋ����[7��6B�!""""�:4¶m�q��-̜����S`�Aa��|��I|��P�j�@�8DDDDD�M� l�:Ǐ'b���P�8���I�� �%%�b֬m�0�#�o#t"""""��͛����o� �3�32%A��V�嗗���۷O����Б�����4��˩5j-�����.D�+=H0��K7��Z�~x�����
Ć�}�U|��^��i4�$�E�~��˩X�~�����CDDDD�5:vl�u��cӦ�����i,�$�}��j�)|��P�l�#t"""""�ӥK�[7�ן×_�&t"��҃�]RRf�ކ�;bذ��i��݃�z�8�Zu
K�:��� S�W�����{����/S`l�ލ�����Y8pS�l�ܹј9���q�4���H<\�P��f�8��(*��W��J��*9**�!�+!�VB�PA&�BM���rTT�@.W<���05���,,L`ee++3��Z�����uS��Zp::i�W^i	�j4�|�g��cʔ�BG"�,=��|��~\����{�sp)�Q*U(((�X\
�X��(EAA���Q\\��cJJ*PYY��gffssSXY���@j5PZZ���
%�˫��{,-M�[[XY������6pr����\]m��d''k�������� DDDD�R�~�QU��[o�ccCL��Y�HD�c�A�"&�:V�>��+G�Eo��P=��.Fzz�����Y���bdf�^��+�R� ������pt����%��`oo	''k��[�����&033���9��aoo##��Z.��V���5(/�Fiie�劊�����V���w�栰���e(,,{��̌�
ggkxz�����ގ��v���#\]mah�U$DDD�l���J��ܹ�ajj�q���HP��A/\bb6���cƴł��C/�\�Dr���b�����"Aj�ii���������������S�����vpq�љ@
�
��e(**�D"CA�����ϗ!?_���bde#'�r� `bbOO{x{�^�x{;�����N��r`)BDDDOlÆ���_�r�(&t"�������vp��O��R##�����2ܾ����ܹ������H �+��d�� W�" ��!0�>>��x���Q�ԐH�u�_����
�G�a��cff�� W�  �AA�?��@��Z�H���H}��q,Yr?�8=z4:� Xz��T�0j�Z��Ip���y_��dU�y3		HH������)���5rGӦ�h��͚y�IO���Y��A$*DJ�ii�	RS�QSS;����AAnxT���qc4h����DDDzn���ؼ��n���� ���;���|��oX��4���9Z$;�W�����t\������```�� W�jՠ�h�ԓ+7�R���U���|��J��HNN	 �����#8�����TӦ���8=��Z�Y���ȑ[سg:��=��DT�Xz�q��m��K�ǈ�Bǡ���A!Ν��K�Rq�J���amm��DD��M� �l�++�@�-�˫q�n�����;��{7II�()�  xzڣI��e���=�����HG)�*L����Eؿ&�����DToXz�s' :z	��i�%K������.$�ܹ�8{�>D���[�}����
@�6h�ԓ�z�    IDATWtPnn	��rq�n��Y,�HIC.W������h��!!�	�Ap�LM���.��Q`����(�޽���a/t$�z�҃��������F���33�`����8q"	ǎ%"!���Ꮞ�c�F	��� zJ.W"%E�;w�q�Vn��Bbb6d�*���qcw�hაo�h�fͼ�{MDD����*���*TVʱs�T��#��҃��3��ĉ$><>>�B��[��
�;wǏ'���;��)���#^z�z�l�6m�aaa*tL�P*����K�Lܼ��[�� �U�����#$�-Zx#,�����BDD�-
�0p�J��Z`��)<��tKzn6l��?܍M�&�k�&B��;��58q"	��ɓwPY)Gx�^z�)^z�7v:"i1�Z���� �-C2!�V��ܤ� i�������r:2�������
�`˖�|�tKz.�]����+1cF��V/�����j�8q����ɓIP(��С!��i���pt�:"�0�J��T	�]���k���޽<(�*���!4�BC}ꇖ-}`i��EDDD�"==��}�6m��v�k��F:��=���2��M�x`��I00�l�I.W����ؽ;G�܆B�B�΍ѧOK��Ռۑ��**jp�F&�]=,C@,.�;-&,�aa~�������q�����͛�6�{���
_=���I'���g�T�0r�dd�ȑ9|���ǋ�{�5��w���h�6���O�V��5:�_��.Ƶk�~=qq�y355
���<,@�-��������]����c�ĉ������c�A�dѢ���g�o�L4o�%t���/Î���X��Jд�'
�����f��VM�7of"66��鈏�����&hժ"#��p?�۳H%""zю����g�¸q텎C�\����ȑۘ0a=�.����Gg(�*�>}?�|'O&���ÆE`��H{��HM�����K��d1и�;���Ꮸ�@�
EDD�l�x���ƺu�ѳgs��=7,=�_IO���//�+����_:�N��+Ŗ-���ϗ��/E��1jT[DG7�������Uaa��E�zU���4ܸQ{J���=ڶB�6�%HÆnBG%""�_|q �֝�ΝS�+t�炥=������
��a߾|A��.]Jņ�q��-88Xb�ȶx��H��M���
\���K�R���8�˫��d��� DE"**���>ODD�/��jL��g�����3���,t$�g�҃����[p�d�y��B��J������xl�pw��""�&tD��!�H�
n��+i�|��))����9ڴ�Gdd ��вe�N=�\�Q�� +���τ���Б��	Kz*?�t}��7OB�.M���u��R���9l�|r��b��h֌C`���J����y�t)W���ʕT��RXX�"<����m�@�n��������O��pt��ΝSaaa*t$���=����3g���9����U��r�f�)��s��0�Ǝmǝ)�^ �� /����T\������ DDDOH$*@߾+�u����Q�Z,=艔�T�gϯѸ�;6m��#i�R��w'p��=4l�ɓ;c��p�A! K""��s�Z��ÆE`Ѣ!B�!�WXz�?R�՘0a=n�����s��`%t$��V�q��]�Xqqq�h�>�'wE���,��4�HT�K�Rp�K""��r��mL���}�7�M�.t���҃��O?��G��ΝS(t��R�q��-,_~��9��=3g�DX��"�W��m�v�X��^ڸ���W�\9
��	�詰���u�V��]�ٳ{b��B��H*�{�^�ʕǑ�,F�>-1c�KNJ��X���/`͚�زe2:th(t�'�҃�RYY5z�Z//{l�����Z��o��Ē%���*A����1�%4l�&t4"zX��>S�՘>}N�H¡C����,t$�'�҃�Ҵi?���{8v�m���
G�;����:�;wrзo+̝��@W�cQ=b	BDD�F.Wb��U��+šC�agǝI����i��X̙��n��ΝGc�?���a�ǋгg3��No{��4�HT�˗Sq�b
K""�Y��e��w���e�d��F�����d1���b����W���������ǩSwѥK����hժ�б�H��]	���Y��v�?���@���X�x��q��KzLU�}�,���)v�OƳ���d����-����Ю]�б�H�!""]r��=��������]��C��Xz�c�{o�c�����A�8��J+�j�)�Ys����7�7��o����`	BDD�n���?7֭��=���b�AuΜ���#�`���۷��q�P���ϗ��ׇ�R�1cFL�ؑ/:��c	��*+kPS�x�sj5PZZYw���&�������f�����Y���.���={fp�i$� �J�Э�b���c��B��ŋ)X�`/����ĉ1kVO��Z���K��dU�H�(((CA�%%(-��TZ{���~,-��\��TZ	�B	��r�5�%ǣ���-``` [[�~������E�es���~|�9[[�=oJ�
�G�EJ��ρ���Б��҃  �goéSI8u�]88X	�^egc��}ؿ?]�6���,i��*A��~��U�033:�V(..Gff�����U���"dg�����UU��>V0��=:,agg�ڕ��ư�0���)LL�`kkC��O���4���a�u�R������XZZ	�Z]�*����n��R�Diid����Q#�UA*�-a��QabggK������..6u�]]m��lgg89Y�N"z"Ri��_++3���4�[D���ĉ$����O@tt��ԛ�*9V�<�U�N����}6ݺ���������Z5@TT ڴ�=��	��))$'���"AZ�ii���*Fyy5 ��������q���=\\l�^�����ť������<���H�UW�T=,Dj/��V������((�A,�>�^�BUwFF�pv����5��j&NN�?ggkxz����v��0���&�
з�
t��+W�biJ����+-�@�.�Aǎ��7���So�K����QRR�ٳ{qni���"\���+W����	��Ѵ�'"#�6m��{ˎ���{7�og!11��"�D" ��["(�AA���u���#�����77��Z���

jˏG+^j/�#EE��ϗA"�"?_��j;;Kxx� nnv�򲇛������_+I��ѕ+i6�{̞��f�: �zo��-8>�O�Swΰ.��*����q��m�?�77[�c=w��2�Ʀ���4\�����\(�*�"22���������Q��TZ����};�og#11���P(Tpu�AӦ^h���
rEÆn<���Hd�K��W�����R��#7���rYYu���̌��a77[xy9�"�ގ��r����֭�!���s�U̚�M�7G ���C�>|&��������u���\��kOcٲ���ǢE�ѡC#�c���
��鈍MÕ+iHHx��<=��{	Ұ���,IV*U�_��x��E�v-))  ����h��͚���6BG�?)+�Fnn	��J��[����ť��.Ann	rrJPTT^w{++3xy9������x���������L"-����a�80���B�!=��CO��[���֭)�.!t����T̛�b���:��0�ޫ��#!�A�)1��"��U���
m�<:�͛{������9��V >^�K�Rp�J:2PVV''k�n� aa~�C�V�zV�����AVV1�����S[�df!'��ٵ�m�k`` WW[x{�׭�c)�����h�4��]D����l�^��Xz�7�؄��t�<�.lmus;��
�}�[�\F������A��u:�FR(THL�ƕ+i�|9��i(**������ЦM ڶD�V`nn�\�L�\�k�2p�|2.]JA|���
4j䎶m�֭}��\�<�Nj������.�;]/((�����	||~?e�ѠZOOxy�^75��D/ZIIz�^Gl�:FF�S��K=t��ML��[�NF�΍���B=z���R��ѿk�#i�Z��d1�\I�+Brrjw�i�ҧn0j�6���y�����\�<��3g�!.N�����]� �k��m�����T��TW+��U�XR�z����Q]���"6Z)� //���q�󑔔��}�c̘v����B�!=��Cϔ�U�S�E��-_=\�8�]~�������	6,�P4"��$+���b���022Dp�ڴ	@x�""����P�=���8>�N%�ԩ���,����vFǎ�о}���|T�/$��Sf��p
MI���|Y�m��M����pu�C�j��b��E��Ɓ70y�F|��H.t�C,=��G���=�p��<88�ֹu;v\ł{acc�ŋ��K�&BG""�ieu�Q��E�u+r���6pv�Fu���EP���0?t���]�Ѭ���K%z��ZQ�*$;�YY�W��ԕ%�V� ���m�JO��w���r��������֬9��{��Eo�㐞a�Gn��B��˰d�!t��F,������$��Z��^XYq�Q}JJ����	��I@zz>LL�`hh��jLM���p_DD ,̏;��V�ϗ=�:��j�G��D��j�G��xx����..�������-<<���l�9��JƏ_�;wrp��[<���K=�T�з�
XX�`׮7u��={��~����/�BG""�*���">|�DFF!���/����022DZZ>��D��KG\����A�R���	�������qcw��#�W]��+@���.�X\�e�X,Eq��[�����E�����bľ�qu������*��nn���)�M��K=��O�`�^?�66t:�3+((üy;q��-��|�
,,L��ED�� &�:bb�#/����!!>���Ri��E�����t\�^�-���BB|к�/BC}Ѻu��s���jrsK K��[R7kD"��}>/�UU��111���5�����jggk8;���Ŧ���l��d��4Vr�}�.ǐ!��AB�!=��C��Rt�������:�3;x�&���	ss,]�*:th(t$""�v�~��-:����B1`@k�>�}+�*$'�'µk�~=��b�Tjxx�� ���	�%n����˓B,.E~����H�((��������� �+���� NNVpv����%���X{<�����%�`gǡ�T������c��>���qH���S�lBB��:�.��M����dUx��_�{w<F���G�{�m����egcϞkػ���Ɂ����o�BѼ�����ʪ��� ׯg�ڵ$$<�X,���!7vG�־�E�VШ�;u�M������ �Hdu�Hqq9���QXX���
��������@�i6�
������ueImQ������G�ڒ%G��7ǰg�t���
�tKw��=���jl�2]�j�n&W��cڴ�Q]-�ҥ��[�`�#霪*9����cq�B2���+-1`@(""����]\�����y3��5��6C˖>�CX�/���8 ��TT�<,@*+Gj?�^��~��zEE����?#\]���p��Z�������L9�w;������V�k��	����c���(*,]z+WG��M�d�p>�%"z���Eؾ=��]Ge�ݺcĈHt���/P
���E|��EHJJ�i1.���Gdd�N1AA�:3��H(�Պ?�!�(*z|�ȣr�Q�RTT�������..�g���"qt����f''+89Y�����\ѫ�d�*��vض�΢����������38{v�ܴo�HT�7�܌�w�����1vl;�#����v�a��X��H���#1hP�־�&�V!..W��?�� ��5pr�FX�""���-�ؘO��^4�\�XR\\�X���2������$e��l �����r���-<<���a77ۇ�����\]mXjj�{��л�2��z'�����$���CGeg�C�/0~_L��I�8Om۶��製p��ߎ։g����R�q��=l�|ǎ%����bȐ�'�yE���Jܺ���x�\IC\\:$lm�ѡC#t��]�4F�NBG%"���>*DrsK!��"'���.7Rdg#/��mML���� ??g��9������h��	��.033�ѓص+3gnņѣG3��b顣�Lل��l�8��.M�_d�*���8��7��w��U���4QAA~��
�l���жm ƌi��_nSS�zA����3g����{�x1�����sF׮MЩSct��VVfB�$��QU%G^^)��J��]���"�D��(Dzz>$Y�m����J���Ф���=��a/�#�?�7o'�#Gނ�/�hz�Xz��x���F���721e�&TTT�oF�S��BG""�Zj��.�b��8t�,,L1th8Ǝm���g�fVW��J�ŉp��]�={�ne��� ��ٳ9��[��7�����HT ���aR{99Y��� ��E�6�@�&�GӦ�h�ȝ;
D.W�_�P*Uطo�V�8I�����Q����w�����/o牨�j���Y|��DE�oF���F�XDDZ���;v\ņ瑜,FX�/ƌi�~�Z�I�?(,,����8y2	Ǐ�Aqq9��=��z5��S���Mii����ݻ�HJ�ARR.��ϫ�ڠ��5�DDD ��}�w+ℒ�U�^���W��X�t��qH����1�w�c�̭8vl.�4�:�?*..ǜ9��ĉ;x�hL���|'"�22
�a�yl�vr�
��a��h��S�hZI�P�ʕ4>|G��BVV1��ЫWsDG7GTT����Z���"ܻ����\ܸ� ��"H$2���Eo���!<��pw׾�ũSw1f�Z|��p�)t�,=tHee:u�ݺc��B��G��ix�͟ �~;��'""�.j�.$cݺs8v,�?�F��������tʭ[Y8r�6��;wr��`���80m�r�E"��Q���ڝ���D�s'
�
����CTT �ti���%K��Nb߾�h��K�8�Xz�eˎb��S�x�89i�v�j�?�p���;7Ɗ#��`%t,""�QYY�_�����p�n.��1aBG��r������[ط�:���}��F������3R(T((��mE�h�Ғ��-L+*j �UA�R���55JTU�Q]�  X[�=�����LM�`oo	;;K��Y<�l;;K�����Ӂ�u�SQQ���u[b�Ʀ���>>��ڵ	�ti�v��֖sA��R�1? ==G��[[�#��c�#��Rt��g��ԩ݄���ʪ��[�����x���x��n|rHD�

ʰa�yl�p���0 ���	͚�0��Dػ�bb��޽<��8�_��0����w��V -M����]3rrJ��[�pG�ȠT��no`` K��[���VV氳�}1cccCCXY�����]��ʪ������GII���P�~:��jOOxz����>>�
rCP�+�������R���8}�N�����00 ���ѩS#t�����;︪���?/{+{��,Aŭ�"�8��9r�LͲ�ae��ʬ�v�rdj���p!�q�ET�%ȼl���q���"p/p���}|>�~���]�~����."t�df�ӫ�7��8�z�$�<B��%��֟�8q�C��hm�������+���.`ɒqt��i���F�βe�믓��2~|&L��^}u���d�m;�?���Ν<<�6�=/��{���@&S������uK��};�[��HI�A�R!�Hpp����%NN���W�;8X��X[[s��7�Ґ���RR�IL�"11���Ĉ�    IDATl���HJ�&>>��� LL�����{<<�i޼NN�|�����.�رDD\���k$'gcmmF�.��bK�w�	������0p����:�@PQ��Q�x1�>}�e������is�֭�x�ݍ��8�l�8� J �D
%��E���P(﯌��VHss�P�TH���B ���ۜ�@���R����#�)���}���O<^T$���a1��HCÇ/�������+�D")[.E__��[C���066��P##�����>z��������!��:��Ո$�g�ƳdI8{�\��Ŋ�S�6�=���6M��;���gٺ�,��Et��ɐ!����W+'=��Rbb�r�F*7o�q�Z�HJ�*󴰷�G�&64nlK�&�4j��}m)�J���M%&�.11w�~�.��i$&f�R���3�eˆ�jUzs����&66���h�ã9~�z��4�_?!���ի���G[شi:~~n�6GPC�G-`ذ_P(�l�<CӦ��L��y�X�����ܹ�������:Dnn��EH��e�ţ���²�Ri���H������g�"�z¯��733BWWr������,Y���8Z�������b̃�),�=��Z`yX@)c|�J��Ru�����D��`aa���ff��oFXXcff����1ss�c��MM�077|��!�JaaWX�$��'oѺuC�N�O_���RR"���h6n<Exx4�����ߚ��;жm�j�'55���Բ�LL*ׯ�-?--Mqs���͖ƍ���zkjjX��V5���\��HT�.\H���x2pu��ukWڷoL�N�xz�{A����g��K��űcB y�N���'os��;XY	1R��ѣ�s�H#F,eǎ��i�is�޽\&O^�ի�,^<�~�Zi�$��Z��df摞�Gj����<��sIK����Ͻ{�ܻ�~<##�!��R��u�&ۥ�z���?f���1�㥏YXch�ߋBcc}���01�{^J����B
U�H��W�L�,K�XPPLAA	yyE����WLNN�����mNNA���"�c����)s�/�WP�_����<^��IY��\�d۶s���n�H�{wo�M��_�l����ز�,6�$::ww;����a��5�Ծ����ƍT�]K�ƍ�2��Aq���ww;����iSGllD�Tff>QQw8�QQ�:u���"��L��w�ϯ	�:y��� r5*�@�����=��n��"�G�3#D��J��_�ﱱ1g��I�6�!Ο�äI+12�g��Ixz:h�$�๑JIJRǈgd䑖&�޽\22��FFF^��� FF��ؘaoo��������[`mm����뛔	��_�N�r%��Edg�E���/!7���*œnYY����զ��1�����!�)h������nW�=��2��F�ݩ�"Vm���6l8�֭g��/�W��Ӊ.]<�}A�T�HH��ƍTbc��o�r����++S�6u���B-rx{;�|0πB��ҥDN��Edd,'O�B*-��Ҕ�	+���i��FӦ
j �
 &&��ߚ�#�hժ����.\H���y�>Z]�A��ѣ�g�%&O^EX�;4m�is�ذ�s�l�sg~�y4��U]�2�����$%e���Irr��mv�-))�0��,��1���{{lmͱ�R�66f�ؘcgg��Y�s	T���rr�"�ݻR�o?Ϟ=���/.�����P�g��咛�pX���66f�٩�oVV����j�������[[3�"���ع�k�Fr��-5�a�(?��X�uQ�L4&F��B��B-t�z�ٙ��逻����xz��u
q��Q(�DG�p�x,���TZD�F6y�M�NnB�<3YY�l�z�u�"��N��ۑ�#�2�]�&�)���!>�l[��N۶���.�n��QCQ*U��|���?�4Z�� ��y��aժ�L�̜9}D��@���. >>������xh?99�\����HggK���\�ԥ����-kel��z�J�X��(��z���F��gڴ�'&x.)��	 ���= ��åJ��J��̉������9NN�
�������ɩ�C��������.�`߾+�pp��D"!-M�L�@GG������ي"�+9s�6׈���ʕdt��s�[��t�ꅷ��,N	jQQwX��۷���HN�>���rG:w���aU*����W����o�qOPn��QC���3̞����
wʌ�<�LYͅ	,^<���[k�$AE�R�������7R����������jMÆָ�Z��7lh-�d	����|~��0+W` &O�Z�+�RiQYΘ��l���%%%���ܲ������������]iyQ3�cgg��C=���� -E�y%QPP�@���eUS���D�R������)%%
��򱳳`���L�X�?�OZZ.�DD\����dg��bE�>����K�6���U�����s����d�7�С�9�c�-��<dgУ�"|}��o�7��\ѣ"�)\H�.|��0M�Ctt2������+WN���I�&	�w��p�R"W�&?�^:�{����Á&Mlqu����RTT��,[v�+c`��+�2aB@Y�MQPPBrr6iiR���)EJ罹��&o��6+�z*��rv����΢F��.

J��+��JB�Z�00�+����r(�6lh]�>^��ªUGټ�::�mτ	���i��	ʃB�$*�{�\&4�"�o��޾�{7�O_����oFPnbc����l�t�������<�+��6�Z9}�6C������0!@��j B����Ys�y�������]]��w��^[[�������"11�K��x1�˗�t)���\$	�ݽ=<�qs���S�/��$'������o����e��nL�P�B���HJ�"99���,RR���&'g��*-������ޢL)�5lhM�V��X��7J���7Ӹr%�˗����&&f���c����:��j]�0P���?�<��#>>�� O&N�BHH�ryܾ}s��5+��u�]K!4�"�v]$::KKShŐ!�4R�XP3����w�ի�r�X,��N��j7l�����ͫ~�1�E���s直h�@���!z�0��dt��9���hԖ_~	g����ё/�xI��*���\Ξ��ܹx.]RYY���Hh�Ė-Т���h��cM�,�!��믇���C�����ݘ4�k���z�&-K\*��
$��ꐚR,-Mi�Њ��qq�*CJ34��v�LAL���cS�.%�L~~1���e�6Jō�M՞���J�T�ʕG8t�:..VL����(hdf�Ӽ�\��t9wn���%�ť�cG�}�7R�J�ggKM�'�!\��Ĳeپ�<��&L���1�j}��J�b��eܹ�ɞ=���+x*B��a��K8����ȹ�JJ���F6o>�G�gʔ@��!�(J�_�˩S�9{6�3gn�������6�/r4�Y3��J.�;<*vL�ȤI]Ņj��Ν�HH�$11���2IH�,˷`ooQ&�<(����Ug�����^M�ҥD�\I����]KA&S`ll���#-Z��������T� �n�cŊ#l�t
�D¨Q~L�ؕ�0��n��n��:��Z�e���ى� �ă%���B:w�`Ĉ����[gV��Gjj+Va��H����R;�L	�ͭ��¥��ѣ�������/c4m�@��G"7��Ϙ0��g�ֈyL�����d�,Kp��F��\rs�8y�QQw8}�6��Ǔ�W���m�6�m�F�oߘ֭]k�ʸ�vQT$cٲ�,Y�D"aʔ@&Obǳ��WLBB�}a���[i�^}}]6��Q#k\]mh�ĖF�l�?�� �)�|9����9��/'��B���ܨLx��Uo���&�TZ�ڵ��\y��4)}����W�ѺuC��i��

�%���tiР>[��^'� j;%%r�f��S��GS��1/��ǘ1��%f	�����M�N�|�!���	�fʔ@�t��y?����//e�5�_���!z� ~�1��Kr��\�\L_�����+�H`���xy9T���G^^1'O�"22���c�t)�BI�&��k׈v�Ӯ]#<=D6{A�B�T�q�)��2���b�N�W5���6���O||qq�ܾ}���t��2���Gzz��'��lI�F6e�H��64jdC�ƶ�
�IJ��ܹ���tw�t)��b9��кuC�7w.�2su�~�
��rtt$���!�)ع�˖���:thB��6l�|��$7�K;9����xn0��IM�a���]Izz.!!>�י�@/Q�B�(�*�®�|�!���Y3g�N����m��c�:����,[v�={f�$ς�"D�Baa	:|ʄ	]�5�W���H�����M�X�rb��T���bN�����DF�r�b
�
OO{:u�S'7���*�L�@P�DD\��O������̚�[�I���E�ť? ��w������A�R!�H��1����RIVV>Ri��:xz:С�ڻ�MW��l+eB��� ��2�ZW�$52�&K�Dp�h�CxJ��������[_�#��L��=�X��ǎ�Ҹ�-�&���166дy��ŋ	,_~����Ӱ�53g�`Р�Z�����J���;w�)�
��=j��z�E��p���՞�q��Ӽ����m�w߽,bK!�+9w.�C��s�p.�A.W���@�Nn������.&��ZAj��?�Lh�E^x�s�����^�f	!..�,OPdd,�o��P(12���X��byYikCC=�4��I��[[���qs��~��U�R(���̦T�h�ܙO>H�N����ڵ�̙�	���zzz��ٙ�u�븸XU�m��s�U���q�i���?�&t	�rq��=��~?[���A+f����!�j���A�_3vlg���isZ�=j 2���?套���/V[�*��ŋ��x�^^{-����+�)�zBq�p^���H�E��X�E�.���ck+��	j*����:���۱�4��/�ҵ�����v�~�.'N����[�<y������u�u놴m�J۶��h��.�֭{ܼ��͛i���q�V��r ��L�Jͺ��n�h�����7o��E�}]]
%={6��Ф�mս!��˕��FrrO�������Ɣ�y�����.A吙����GY����2�kϫ�v�Q#M�&��ť����ټ��Ζe�GM�����3̜�����&��!D��g޼m�:�Q�)�
��9s�fÆ�,X��G��@u�����X�ơC׉�K��ԐΝ=��[��4n\���&HJ�⭷�$2�&�'w��w_.�D.Wr�bB��q��-����0�}��t��FǎMh�ҥB��J����ln�J���{ܸq���4bb�.�kbbP&�xz�//uiZ==v���)���%���.J��ѣ;��;/Ti��m�>����8��t��Rb�\�(,,a���,]Abb}��2sfO��5m��p�N�����ѱ>o��С�k����kp�x,���bi)��j�����Jгgs��X-}�d
f�X���WX�l=z4��~��͛i��]�����<y�B����5�m�F5�OQ ({�^f֬���3��o_�U���6��QT$���;DF�r��mΜ�MAA	66ft�膟_:vt��۱ʓ���p�F*11��Ʀr��ZIL�B�R���������e�m���.��z��FS�bd�_�}���w˼L�==]��7�ިOA�P(	��?���/�2kV/!~�EBB&?��ƍ�pp�ǌ�1�c��ΓJ��c>>N�Z5I���!zh9�7�a֬�8y�jɰ^XX¤I�8{6�U�&U{��@s�d
��������]%..���M
jJHH3�D�G���$11Q�fh���_{=�d2���_=̰a�Y�`���&���>}��Goy���;�d
4���O��ѱ��Ve�/((!66�L	�������K�]]ll�������/;w�@�x�P�ܼ)���l��K�J���(F*�ST$/{�D"AGG�D�B�P���̞�KÆ"GDe��燋�K���R�س�2�����d��⇠�$&f��Oa���I��,�1�;#G��8�������>��c;i�� D-F�T�%~~n|���*�O*-b���ܺ�������[��͒��Ǿ}�	��С������H��>t��C�v�j]Y�ʤ�縩���������d��r(��մI��\Ʌw8z�G��p�L��r�4��S'w:vl���;NN�5mj����s�����\�DR�[���LqqBU��D����)�������7CG�}}[������AQ��*���1a�V�\Ym��T*���7��O�x��xz:T���Krr6?�ƺu'pv�dΜ>��תF]�,Z��%K"ػW���C�ٵ�Ӧ��ȑpu���byyŌ����L6n�.�ZLRR�w_b�:u}}]:wv�G��{Ӡ�(]X^$	�֭c�ȑ�6�ZY�~=�F��������5j9 ��>YTf�T*��);v�7G,yy�88�# ��.]<��٣F�RR"���]���}��H��ӥ�D�}!���޽?��DA53j�( ֭[W�}�����ڵ����ٽD�bA�HJ�b��P�n=K˖.|�a���P(8�G��d���U�U���=���T*~�!��T��QPP1˹s'�͛g��&���͛i��}��Ћ\�����!!!>,]:�� oLL�۾@p��mƍ�77[V��,�,W"�o����;v�c�b�����ʔN�����~x֚<7o����Q*n�d
T*��:4jd���>>Nxz:p��if������H$��݂�=��m�y��2��9Ǆ	]x���
�e���-���Q��j7,��K/�Lp�7s���iS������_��5��Oh�$����~�+W����U�Oa�Z�y3���~M��˗��Ȟ=��v-kk3z�j��o�& �S(��=øq+���GUIbɺDvv�_'"�G�� ))SSC���x��x��턎N�q�./���e���:��XѼ�3^^�xy9���@�ƶ��=:��u	�}�S�@GG Amx�Ŗ�Ys�o��Ǻu'�1�;�'wc��4o�����r�H�~�����:�=o��[���\\��⋗x��u5���0B��R�,	�|�Ե������W�ʦM�E�gG�Tq�\�v�������-�ի9�>����c8t�:'��_��|���;� 
����;��Gs�pQQw�H�]�ƌ�G�.�n����~m�kW/��zm�6*��"h���L�ԕ#:�dI����?Ƈ�Ȁ�kT�A��ɞ=�پ�<_|����/�81�7����X��=�����̙뉈xOx7�Q�衅\��������f��Q\,g�ĕ\��ĦMӵ�EM�x�r%�����u��{/��*�I[^|�}��Ҳ������ѣ7?�7j��_��3���MD�5����1dg��bEPPS�O�sg,,�4mf�ch�ǨQ�����v`jj��o�f̘N|�e(3f�eŊ�̛7��m]5m�@��ё0p`��mɪUG����_�7���ĉ]00о��C��9s6�t�8M�#� ����믇h�ֵ��td2�&�$**�M�����T��v����Q%6	*�ٳ�bjZ��u�[bj�ąQ\�P���3�~��U~�u��4Tw�U�wM���;L�����۱h�0!���rN��ɡC�8t�:��)Щ��g�"0��H�]�<�����R�گ
������[�x�&N`޼���{j�G����B��	�}}]�L	dĈ��s8_}ʊ��3���ժ�Ec��n$Ç/�W�s�F�&	�!zh��R���?�X5�<d2�'��̙�l�0��͝�}�_�ŦM�:����
�G�&��12�Wy_�6mB___�ρ&/�ń�a���;�W����ꫡB�x����_%<<���oRXX���#ݺ5����熡����i<(B�A���)���i�ܙ��~�ݻ/1�6�tY��ݙ6-H+W�ڃ��1�ߗ	���W�y��?Y����U^C�t�m    IDAT]�x0iR |�?�&8:��
a��!F1-c��#��YЧ�o���R�x�?9y�&��O�eK�gnc�ȑ)�&�<�%����TZ�ȑ�pu�fɒ1"���r%�O��������7R��0�[��|�� ����E����-
jʲe��l�x��(@
���C=/�ԩ��������=Çw`��~XY�j�< >��E��[o�ş�*<�B��"�����c��f�*I����ر#�u�^�M�Q^Ms�Z
��7	
jJ�F6U�ϣ+���>�J���8W�ǭ�V�K�6�T�x�5 �_?ccQ�933���h�����אJqw��g��|��Kt�ФN$ ����o�����}pyt|(�I�g�x���1�q���q����*�x��v�f߳�����ŋ	=fjj������>�����a�$�52�g��ڞO>���_^J�~��7o�=�����6�ƶm�?��y�>��I�FF����(����U��2qb�F�TB��"6l8��1�� ��ߏ�������(�t��������GY��8 M��ҧ�/�z5�uk�*�I���W^�����^,^���ț���f�L�YJtt2aaWٿ�*��ǣ�������ݻ���j�i��YˏNڟv~e�S���>˘Uz�IB���K*�<�ի���{�3�Wtuu03S�g�����>����!z��al������`h����>ffF�ajj���!ff���annĢE�1�}���]2{vo&O�*�P�2`@kBB|���}̛��y��Ю]c��ղ�3g����w腛��EU����T���Ì凩�a���o�e�������e�ඕڶ@P��0F__�Lέ[�X��?�t�����ݻ%={��U�^=������Av��w��c��qu�bUQ���Gov����$'gcggNHH3�M�kW�J��T��[�H_z�Tv�5nVǹ���|��w�#���y��%��'+F&S�P(��+ /��BAI���� rs))Q��_LFF��
��D��eɐJ�()���_�D;���H��O���סxy9��b�����fXZ�biir�f���)���kzu_�9LM�;���0�-�##G�����17����o��������:�m�)D�:�=��������Y�nV���3m���ό�+�m���`ffă��%%�İ�مl�|�N���K@�'�{��G�fϝ��щ�������Ʀ��[�6-�_l�is����|�®�w�e""�Q\,��ׅ�#�	�E�"�Y�/��;�>j��fh��T�������WDn����SH^^Ri		���s����)�ѱ/&��U@VV~��� ���++S��Ͱ�6���66f�ښcgg���vv��{6l�����;w�|��p���j�==~�q4=z,����3{v/��!�>��%���!�����ٲ��LI��WV��g���v�G]
;�$FF�O<&�)�o<x�C����{�h���z�z�PTΊ�|֕�j]��J��8q�[�2gNM�S�ܹ���}Wػ�'N�BOO�.]<�?`��u��Ou�'O�C�o����SSç���ٴ���o��D�_�DH��.m���Of�ZQ�
��T�gf�s�n.�!##���<���}�FF�	!���pp���S}��-qt���S}QQ��ҿk:w����0z�r����y5nڤ�-s�ȼy���ݛV�V���C�Z���I?ˎoVZ�Ri�G/���BT'�:�J����(*�#��w�-&?���Ria��nn��u7/����d2�����),�����R�,G���H$�����I3��ez����I@]�L���_�d
~��v���.%�o�ev��ի�ԫgB���������E؊��T�8���Bui��
$	Æ�'8؛O>��ر�2`@k>�t066f����޾^��R(�dd䓑�KJJyܻ�KZ����<�_�����IIɦ�X^v���9���qp����%NN�qt���s}\]��ݿ����6c�ұК9s6q��5��z8ݻ{W�-��wa��+̜���{g?uLP�����o�h�ֵ�jY��J&O^Ivv!;wN�	ՎLV*@�PR"�/@���"�)���999���rs�����QX(���,>9?����
c�011���CCu7##}���qq��ܐ��BC/�g�����d
���?�c�ba��B�[�J���+��o�v옉��v��{^�r%'NĲg�e��LRR�Ζ��ٜy����.��O*�K�*Ɨg����XQ�>m�6��T666f����iǜ9�\ȂC0�u��������;;s��������<RR�II�&11��d����I��w��T)2�:����>���4lh����#�6�)��y����1w�ƌY�С������$�H�	
��v��7���T/��a��ؾ=�o�Qim~��v���m�L�(-V��o���y�R��<6���'��_��ڞ�GE�y��<�D��mS^}�wJJ���b�����=�u�_m��H077�/@�aaa|�,�ڭ��@WWk������z��bb��L_��	���������<����ݗع3��$	��jȐv�Ӊ�͝3�ټ<*�t���)O��;��_̟?����駃iѢ���y.��d<x�]�.v���||�6�=�{���OP1*���icCyǗ籭"��cge����@p�7����;�>�v�b�¡�ؘUj?66f�ؘ=q�S�T��I��� >>�;w��ر#��Ti�s�����jM�Fָ��Ѥ�-��4jdS%e���~}~�i4�����6ҳ�"~�ym�T�Bpypp��g�b�����bK:thRm}�!zh�NajjXi���o?ϯ�fٲqx{k�:AE�k>�y�d�2lZ�*�<�{P��*������]�J���ښcbbp����}�� ����xjQ� SS#�[�~�;���.r�__gƍ�B�~�D�@";��W_]͋/�d��N�6�B��~�]�.r��U��d�oߘY�zҫWs6������n`jjȂ/ѧOK�~{ݺ-d����߿U�� �H�Bk7q-*��D�FN�:IBB&
�==6����ww{������aaa\m���ѫWsڶměo�g��x���1�;::Փl{Ȑvl�śo�IX�;��/�چ=4�J�b͚��r�JQ���Sx뭿�6-��T'��2��z8<Kϻ*�<}?x~E�yR��+yyI�����Ն6bj��s���`dd���=ڿ��ç}�b��|�T*f�\���>_}5L��<99��{��Ћ:t�B���;<�޽[`gg�i1N	�H�.����g�mgڴ5���_���u�z}T##}����r��1�L�͛i�Ʀq�f11w9r$�U���U���3���{||���q�iSG1A�$ll���W���|��N���F��P=�Y��z8ݺ-d��]"̥"Dr�H�������Ri�&��}�Ƽ�~�J���h���\J�6���Hi���ӧӿ+�%��t���/��s��BCߪ�9��y��s�]�.p�x,���]=Y�p(={6�5�H���>��33C.J߾-�=�/�w��o�����A__��Mi���IIY�!11�l�r��	��Ь�Z)�Uf5ƺ�D"�W��wg��5t��5�~;��=�Wy�vv�|��:̥O_��ܪ�OA�!D����������Q�T����r?�<Z�Tvނ�@m~m5+�][ \Wk�]g��P/���<m!55�]�.�k�N��������|��HBB|�5��@ T�8�.|��ѣ�3iR ~د�%uv���ْ�@��OJ�����ۦM���KG�TaaaL���x{;Ѭ���.xz:h]x��Ҽ�3{��棏�2a�J&N���Wy��!Cڱs�f��K���2j֨S��{7�����b���nk��;�?����OCe:+^R���ʰ��~4��k*B����g0m�ƍ��С�5mοHK�e׮(v���S�055$$ć�K��-*m	�Z���?�8��`o�ǎ�য়�hE޹�T�ѣY�c%\��r_I�ҥD6n<Enn&&�hр֭Ҫ�+mڸҠ��y&&|��p�x��t)�e��aooQ��~��0�R���X�.�zt���\턅]e��},^<__�J���h鷚T2�Ym}�r}�ӏ@P�(((a��xy9��'4mNy��y��;�8q������ٜ�+'ҭ[�g�4$5�A��о}c^}-}�,f��~L�P��}MLh�����#J���7�8�QQ�DF�dŊ#�d
lm�iժ!�[7�ukWZ�n(a��V��81q�
z���e��Ui���0�7�X�/���/�\j�jK��J֮=�ĉ]�++qbb�����c;1|x�J��r�h���>�Yx�>��L^e��+�MU�>	ڀB�d��?��.dÆ�/7���Oh�E�o����X��ѣ˗�'(������&i�����~�c��m��G��#k}�fIY�a��^���r._N���;�?�ƍ����H$�4��m[W:vl�����j�hww;BCg��[2t�/|�Q&O�Ze�Ҏ�Ћ̞-�\jB�� {�^"33��_��p
���3���j-\�A�f��-�8�֭o`c�����v�ĎQ=z]]BB|X�d,ݻ���@  �����7{ؔ�^���ݿb������h۶m�6*{,++��7�N���Gm���{{:vt���7<=�k��Ly033d��q,Y����8w.�E��W� ��C�^��g���>Շ=4���O��8���p.\H`Ϟ�_��fJ��j���ŨQ�5j��ͨ��Xq��k#Y�rb�ǈ���w�e�m;�����ё��?�"$ħFT�h&&&��W��Ht��1F"1@G��������ꭎ�1�����1$3s��w*�~==K,-�����< }}llF������R��4��}���).�C&K�w�0a�5��ѺuC����s�0~�
Ǝ���������)���{j��8y�&'O�b��]H��XY�ҡC���B�����1�*$	ӧ���´ik���{V����E!���9�>�3�ҷoK�RÑ���Z��K�s�l��Z�K!EE�a�����!��_�>�҉ݺu몭O�� >�Ibb����4�߿�ƟǱa�)f����0n\�j�S&Sp�p[��eϞK�d
�ukʀ��ѣ���"�0r���۷�P(�鼹sO��+{�1�D�DBY�J�B�T��ߧ������&�
����dv�`���4ibAvv1�|r���k����s��(*6m�Ett6��Ř����c��w}�6����ɋP~~~��h_�5m`�����Flm���14k�i���REtt2'N�$2R-�dd�ann���]�x䍻���M�����8q%��Y�Z5�!���dҤ�DG�p��;uZ���ѣ����Pv���#�W����bz�XDӦ��\���_�1�ۈ�_�Ml��k���;��o�Ti_*���g�غ�۷G���O���4������ҴJ��ƈK8|8��������Ǒ?������+W�x��u�Ĥ�T*��4�ҥ���+�_�o�q#�ӧ?�ٹvU��r%���h�ã9s&�ڵkLH�AA޵�:Iu����믯�ܹx���%��U�-�T*n�H�ĉ[?������.��Ŋ���t��E�.�XX�^1����7�\���WX�h8C����>RS�t��%/�܁�?֞D�gC��T#J���O3aB�
�1w�
K���h�@ ����믯eڴ�*<n�He��sl�z�����x�@n+�
�����]n�CWW�Ν�Y�b�s�����۽���$�J%�����B���q�vF����j_�W�f�4k��믇��]����	�ʒ%|�����	 �"���X���pa(�f�ŉ7Y�`�XY
�OO<=;�
����;DD\�С�[w�L�+AZ�h�\E��-Ǘ_�2s�zbc�x��*5牽��|ҟw��H���iժa��-�>��G5r��5Ǝ��ӧ?�P��;/�꫿�a�T�t���X�ۈ�_����9f�\�ر�����O✚��֭�ٲ��/'��X�A��0xp[||�*�?��2
��7RQ*�|I��#aȐv,Z4��r��:u��3ד���B�|��֭3�������\��c���L�1�R�ŋ	�����k\�����.~~n{ӣG35�Ѵ�ZMX�Uf�\�����6AT/� �b\D�5�!%%kk3��&(�i��Tܼ��go�g�f��èJ���R�1b)��"�bE���ԩk(((f͚W�����l�w���#;��G�����FLz�6��h�u�"�3�o^}�s����v��"BC/�e�Y����ܘ�}}<�-~~n�jULP�(*�1g�&����E���|з�+����,X��ի���#���ammƈY�$�!;��t�sgQ������MDD4^C*-�Q#z�hFp�7~~n
��GIJ�b��Uܺu�E��ӯ_+M�T㉎N)��:u�R���;�{��O����Ӵ��͙3��8q%NN��Y�J��C��Ϡ{��x���V�JkWP=ѣ���.�U�O��1����L�T*�_JVV>��oiL]5j�6mҺI�\�N�f`P72W?YY�XZV��xԨQ:T�>A�`�҃|��v�}�f����핔�9p �͛�v�BB�1dH[���10��v���5�X��$��%H$갓�Q'4���ȤI]+����ט5�/������hU__�����
h��F\��E���M��JΜ�MX�U""���N��Ā� O���		��ɩ����JJ�̟��U��0aB ��+�D^^1��W	�Hxx4��%�iӐ޽[зo��t�N�ǯ����u�^�I���Z���d߾�xz:TZ���G��ĪUGY�x/���{�{��|��f���*��;w.�����/E"�C_�g\04t�����iӴ�� ��(�SROqqJea�������Ϫ�J��ad2|����:����81��m)�*"#o�e�Yv�@~~1���Җ^������RšC�Y�����88�c��Ό���?`Ŋ#�djQB"���#��Gӿ�
���]�'�leӦ3��sw<	�c=M��-8~~����$'g�	 ��PXX���c� Ү]c��ĂΎQ̞�^^,]:��%��4��r��!4�"��]&33��M��Ǘ޽[мyͫ���S��	+�q#���L�6��ҮB�d���H$l�����Aѣ���s���̟?��KM�!0�K�N�ƛo�MW���bΜ����[9r������]�-\8��c;i�R�4�աC�9x�:QQ�(�*Z�h@׮^zѾ}c��"����2e5����_�УG�
�s�J[��e��sܽ�C�<�-��ڏTZȆ�X��qq�t�����]�ի9���I����T*tuu04�c��Iϕl�ĕ��s�ϔ���cE77[����6����8q��v���t,,���M�{!8�[��sկi�Ʀ1e�jRS�|��HBB|4mR�D�Pr��-BC/�w�e���h�К>}Z0hP[Z�h�i�Mq��3��ҥ�*�;s�Z
�z}���.:A�"D�j���dBB����w���٤I+���`ϞYuf2��S��S�9q�&G����B�zH�(EWW�)S5��&#�q��T'���K���?�&t�֔���u�ֻ@���Mcܸ�()��f�d���-�hjj�}�M��s�F�l4����kA�!::�ի��y�D�&ty�[��!?���	6L�Y��[��~�.�ǯ ))�Ĥ��y��d˖.��=�쨋�ť���ã9q�&2�__���ңG3|}]��*saa	|���O3{v/�z�g�V�<�J��v�ĎQ�ť����K/�cР�5"K�P���������a�ѱR���=,]z���wqq���6U�=���>���ӷٳ����w��ԩkرcf�(�TPPB��G���W    IDATff> ��@���G�����.�Z5d˖e+]�����C�9r$�#G�#���X��@/�uS�z���=Y��˦M�����4m�Ȋ˝���D�޽�ٸ�^��܈A��2xpڴqǂ�L�`��K���Q"#o��n���]:�=��O�:q�&��7�WO��պR�)((��7�m�9*r��Ɇ�*Ŗ�JAA	G��MX�U���U8����C׮^ԯo�i3���k#���̈́�����05�}%����g�ؼ���s���N��2�}������?�Ɨ_�2{v�JIBZR"�W�opp�ǟN�U�=��LA�V���;/0~|�r���S@`�Bn���B��\IÆ���\,-M8p��J��,P#Ba���U�W^�ʇ�+�w���86l8������/�[7/��@�^�EBRA�!--��k��vm$���ңG3Ə�L@��Vvｷ���O <T�E�����^|�%˗��b����)��_���hΜ��J��5"8؛��}�Dy�ӧo3y�*���X�rb�N�Y�()�q�M�Nv	/�Ђ���ѭ���.Dn�p�w��Ș1����A�=��=���?�x��m_IV
�
!zT1�v]`ƌ�DEͧ^���f�ŉ7	{�*�P�8v,�a�~y��l)��:l��:4�&��6O�	lJ�n"F�|\�������*��^�����+6�"66ooG^z�=��y:5�3gn�b�BC/bnn�ȑ~��I�\�cb����ѭ�7�O�"33�L���.���ťSTT�J�p����C����o_֠����������Fxx4�����X�,�K�Z�	������+HH�d�ұt��i����������̙8ll�4��ٻ븨�.��@��V,�VBL�������5^um��,�.PAlQ$,D�@@``����]W���~>~֗���û,�ι�9���5NuYjfpv�e��=��рի��;A3�IN������:�I�6b�5�l�>4��qs{̀۱�K�io@�]͜y�#Gn'Y?,�HX��;�G���Ȅ�D)��,��r�mse�'��/���C��̟T�J�~��խ�ɑB�EE�8y�w||ޠ�WK�t�n@޼YkwRXX��k)Q�G�����(Ǝ݋�� N����ny��9���ބ�}K����.e���,Y�K��E� �+��zťK�8;����
55)M�V�]�:�m[;�=����1c�!Μ�d�<3ƌi���aaQԪ��z�y�`��K�p�ǎ�%  �F�*3d�ݺ�g�]���6̊���iӠt�Z����e�WgÆ�J�RP6���@aa����۶�s��)zϷo1�k�M�Ve���a����G:w^˗/�?u�WWW�Ĥ�vSMp�OD)��V~~AL�fǣGA̚ՙѣ[':��������I�~��+B���e({�^�����1���cii��q�ʦP(6�
o��8:�H('��,]j�޽�y�x9R������n�r�ْ�{�s��]��dL�؎9s���;ɝBC�qu���E?�^}��ϑT�T�6mjӡC�5���li�u�+˗�Mx��7�:2Y��m���g 8;�Lws_!y
��kמ��u�)T(��7a�#��J��w_0x�.7��Ν�ȗO#�k99�0|�5��M״,!c��G���ɢEg���3�7��u�np���*��)n�xƄ	��QC��W�𚺺���YY�aRn&Ja�����ٴɅ��/��[�u���3���+ժ��_�Ƙ�7�+B�"�+�z���n���Q�ta,,�3p`SJ�(���~i�G6nt�ĉ�VJ��ןbn��fR�^��ʰ�(Ο��ظz�����'�Ν\���ŋy��-��yh޼��ץM�ZY��*-._�gܸ�T�T++K�,q�����X9��R��u8sf����U���8x�&� 8����e�4jTYա����S��6{��L�g�#��������H�iD�#��
��fM���e(�Z�`�ʾ�훻����Y��68ӡC]֮����Gpt�&6V�D"!o^u��fP�ziU�+��(��������1�?��o��2jT�������t�n��y�_~���(,���fϞk�`dTK����˲�����ٗaìX���7�屖�V|�űc2):!���>'����?!""��5�i׮�[עiӪ����B6�
�,�����􈓰c�P���U_n'��ћ;�p��6�̸qm01�����O���_�m�)S��Ǡ����u��>Ӫ�
F�l��ٝ���"�A���`h��C��al\=E�>ܚ�8sfJ��ԞY޾�̄	���|ɂ=�܄��cd����( �oJ�n�UH��,����++V�cԨ�ԪU&�����/>Ñ#whѢ˖��J���(_r?� ��q���H�z�n���15jh�:�{����k��E?�7!/c��a���fR��2�dqܸ�4��ٳ�hi�E���o_�6mjg�Iy�d֬#?5ŗJ�dI-nޜ/�ƫ�ݻ/ؼ�_*W.�ر��۷��ʠ_��O��-Z�#Gƥ9�am�ƢE�qv���~��"�Av������X���ի�8pg�NCO/�4�st�fƌ�/^�;,~��|���L9��e�.��re��;v�ɓm�7ό�cۨ��O.Wp���/?K��yX��;ff���Eq�����(_�5�,GGo��q�ƍgT�Z
KKc��iD�B�T^���Gӵ�z
�éS��� 2o�	��|�qc^�� �,  �K��pv~ȍO����^�r�o�U__'��V�y�}�l�a�򿩩I�>݄i�:frd�={���[/q��]J�*�����O5ɏׯ?ѻ�f�-���c��b .NN�nȓG�'&��فHzd�N��ҬYU,�챱�r:v\M�Y�:e�0�]LL,��fϞk��߄%Kz����hއ�R�zi�3HO)̄	�9sƓ���r(��l�:���4+7�{�������F�b�t���bk{�3g<��M�A��Ұ���{!�޿������·_i߾��ƴhQ#[��*
F��˭[�pr�A�2E~y|DD4�6̈́q��dR�Bf��-�kמ���˥K��z����ҪUMڵ�C�6�(R$�߾����l��>m!t���$� y�s���d�����M�\�����va&Mj�����ן07�B�92.M��7���e�rs�uY���D�#<{��-���8=Ec�����_�\�6��ųvS3ec�H?~ǪU}��]��?KM)�B��n�y|���~uu544�,^܋����;�}BX����{cdT���½{�<x�Ǐ�Q�~ylJϞ�hie���� �	=kkwΞ}@�B�0�)C�e�F��6��z�#���iӪ�om����g��X��-�B�������.�q��s
��סcǺ�iS��u˦(�d�=[��R�\Qv����N�c��q5>>o�=NCCSS]�m��s
����g6nt����څ�6�#��2uٿ��KSBo��3<x7�?�|���D$=2��Վ�>}7�?�=644��͗1c�	�F�ʄ�T������hjj�g�H1�CH�_��ԬY��[]zO����֭k�~�@J��>5��QX�7֯�����+��ܼ!���9/��U�{wn��d� d5QQ2N������7��U`�0cz�h�#�\��ϐ!�X��;#G�L�x�\���2ڶ�͒%��47
����..�tɏ��R�taڵ�M�6�hժV��8:uZ������P̜ٙ�ۥ�l���Wl�|''@A\���>�H$N��$vfAo�|b�F��nR�J)���Bǎ�2����[��J[�#22�֭WШQe�l�AQ
�%���h)���>�$�cg�<���Ϲxqv�/�8u�ӧ�iӪl�6$W����ߥ0/�� 66.�c54����Ú5���E/�#����d�ظ�a�3R��&M���D``���4�)ff�( FM��˗���{�C�n���>���4hPQա)͋��y-&&�ٰa`��������ָ��A��%38B!�S(������!��~ܿ����&M�ЦMm:t���+$$=����hT*�/Kݶm(�˧o��O=z��{�������~�?PW�R��6NN3E��,*  ��K8w΋&M�0w�����{�{�P�|;61ջR]\2t�.G�52(J!5D�C���I�.�~}.�*����ޯ��y-��chժf&E���r+V�e�WF�j���ݲl,!{��k���l��u&�HP(��i���梬B	d�8�źu��)���J��y�ݻ!6�vm1IG�~
W�<��Ɲ�R�ta,,�3p`��]9,,��]ס��ɉS<1��|y�s����PȎBCùr%~����|�I�
�h߾.��l�~	���k����Y�Oi�����3g<���	�J%�Yӟ~�+�\B���d�2{n�|���.s�vM�3�2�y�=6���šC�R��f�k=z���l1�.I%[���n=�����ۿ�v455���	��Fxx4&��ʕG�\�G\X����Q���d����/uu5��ϦM�E�=��r'Nx�r�9��>�������6� A���E/Gl�r���(�Ş=�O��7���e:v��#'���ɱ�������MC[;e�����h�v��u�Z���}��u�/�.����7����v z�2dٲ�J�~ř3�ٳǝ�ߢ���L�T*��oY����9;��t�/^|`ܸ6L��>�w��г�f�U+ɾ}�����7o>Ѻ�J&Nlǔ)20J!%D�C�
M�.a�P#&Lh��c�ݟ0`�v.^��cg9�z��!Cv��K$�w[bhXI�!	9�����#M�-W.�ʕ�(9����-޾-�B!A]]N��hkG����u�����������b�w���D"�ܼ!���9���ݲe��y�'&��\g֬#ܹ�K�fg�)5����ɩUkѿ<N]]J�RZ��a��a%޽{Ǵiӈ�K��_����ݻ�O�+_>�J�rƽ����֭C[;g���g�;�W;��������ٳA��z����[�ӫ��͈T�#غՕի�|�71MP�r�cz���^}��T���)����s����ۿgU�q��4��2��� ~]�<�I�NI� �CS3-��R����KH\�r�뿧v�4nD��a�Nx=z�C�))BAH�L���z��L�v��~�)s�t�޽�,_n�c��ߝ>}�-[\Y��o�?Fp��]F�j)B�yx$�������a�豑�k�pv���kD�2�V����[j��D�RJY7+8t���?7v�)�ե�ْ���ҡC]&O��[�xy�ʰs֬����X��}�ر{9��F�jEŊř7�D��'����Dg�zQ�n�dz9:�����;,2)��u��SF��FW���Õ6]cbRw�'�n]�"E
P�h~
֤H��)���E�S�H�������V��4h��Cr���r����·_i߾���E���C���k�O?ĨQ-�۷Q�޻o�545�лw��N��\\�'�:11�'ʿ�\�� 5�B9r$C���r��b�
�jU_�m���'05]���1��f�!=���+���X���ɶl�8(E�	54�X��s�-8:zөS}��&��Hz(�ٳ����7qqrV�<ǰaƔ+����Yѹs^���Ν�q�?�FP�F�*��|Ar��w_`c㎃�
�G��M��hN�
�TZ�
g�0+5�����R�^�,��{�ѿc���Ƞ��l۶K���QWWC*��d<�WTRؾSSKY�!��W�'NL�ر����Ν{��E=��M_��24�Ȟ=#2d��`�r���Y����m���'iٲ&��/��<"�$��o�k�_��<v�.AA��4�}&E�yN��ǤI�f̟��5�fA!k���q�{�\���5zzX��/=z4ȕ�ve�8F��!o^uv���Ij'Nx��c�F�ʠ���K=BC�R�RI
����|,�--M
��{�߿��B�49tȎA�֫:|!�H$��ӈ���d�����ȑ�,]ڛ���G�Ȩ۶a��/�̙�R�����;���X��s�vUjLB��+~9{֋5��^�t��DG���_�3�5Ŋ���2�ѣw�>�cǶ�1� *��e({�^�С�DDDcf�ϲe���wEN��������S(\8�ޫP(ض�=z4H�A���ۇ�:!�*Z� k���_�F���1ڴYɬY�5��R�ou�X�5k�3m�%K�¢y��)Q� ��ޅNҧO��阕����88xҭۯg����NLL,�G�Μ�2���Mf�:����=����Ar!�B���c���qq�t�Ӛ�P�d!U��r66n:tk��Ԭ��n��<y�Ν9�� 9C��Upr���m�X����YӟZ��(�}�6���0��;���&={6H�=C�4���[̙s��Gǋ�LLoQ�Ǐ�����_Nm���f�&&O{?~��3�0}��Hx�ʯ.V�B&�'<<wZ�ZA��ۉ��b��aܺ5�ɓۋ��S�.<ͬY��ر^��ر�2m��O(�\G"�$�'-k���B���Pc���8;�D*�`b���k����?�����1vl�N=�0I�W�Ԥ�Xч�7�ao充8��;=�����+��N��I�w�5����СF�Y�:ޛ�S�0�-ӧ��:A�2
E�׈o��u�%��#ϟ��ڍ�G�'�w���9L�O�r���ƍ�G����<9m��<<�~�)ǎMPrt���$v�K�����⿏���U�ziN�����WY��g�z�a�@��+������Bp�,,vs���d���U��&,^lO�u��MM3���g�zѥKһ<��d��q�	ڑ'O��3]���ر{:�9s�� BƓ�\��À�i�b9��~L�n½{Y���Hx�GXXC��b��[7 �O�w츄��FFՔ� BƒJ%�݊�gQ�h~�tYǺu����{m�DºuhѢ�y��S����.��}c���>��r"�N/^|���-]�$=����R�����dbd���5#F�Ы�!K��Tu8�����ʚ�k����H�o�Mo�����xRsNAH�/_"ٶ�FFK���F"��w�H���0fLk��4Ub�+g�Hk"#c���L�ŀ�Ν�b̘6J�P2��J{-��ߤ���?Ss=�Q�T�G��g�<36mr�G��<{�>�목Iٶm�Jiaa�����__�xA�M3a�VW^�M����I�trr�E[�0���}]&�c��K��&G��
�̰aVVdժ�◱��}߆��Ob7%I���5�z���הn�Mi�ʌ'5�����{ˬYGh�`��_�}�:������ch߾R��%e��xx��(J�N�����/��S��]�~�#Yѯ�ѩ��&��#%׸��ߵ�u4�I$F�jŅ3���ӱ���������f����9�:��!#F��B�b,\x:]�RN$=�����zI~�9t�11��,�#S���(�I�"���=5U�$*��e���Z�<���r��X9��{3���ŭ[Ϙ7���,Yҋ*UJ�:�,���*�`۶!��7����r��F�n-LB���kҿ��=�Pq�8ժ���~*�Ƿe��S���￦k�2e�p��h��^1m��/��ih��xq/��r�Q��+��Hz���ϑܾ��v��$�zl��-[\=�U�oT'g}|������ʧ�!�Hk������A����l��B�&�;v/�
ir��X�\�KK�5�,#]������7�4Oj�n׮+hi���J�N���p��
1�V��Rf�0��~*/_~�C��ҝ��]��vYr��}�lq�屭ZդS��,XpJ)�E�_I�t�tɟ|�406����'Oz��s$Ægrdʷf�W�>��j8e�Qu8�����鐪%���
Bfx��S���p۶]�G�_�˞=#hٲ��0�
~~AL��s�L��.]k��}c߾k�Պ|�4�� dY�ڜb����*��4��-k2p��.uH�h�-j�dI/�/?ˉ�<v�����w�{��'���    IDAT�L�o2�B��޴hQ#ћ�\�ƍ.�ՒB������g�a�3k��Kv� ���]e��f���4��$����� k�xxR�vY�.�E�^��~g�����ciiE�z�Y��o�׳�qG"�`a���Br״��?#+Đ[,��M�al\�y�Np��S�l��N�4�gaќ7o>1m��Ji%��\G�8cǶ᯿�ѣŋLϷ!����F2YW��Ӿ}�-�-392�z��Ӧ�1t�Q��>#do{�\��h)�����;x{�&::6C���f7��e)ih��5R��2�LK<�%BRsNA�.88�իi�hS��R�L���ŋ�4��Hx��LǰaVH�v�Hwϭo�bص�
#F�eEB���kZj���52��z��O\G��~�s��t��b��q���i^�?�е��F�!  $��&NlG��yX��l��%$O��H�[���d����.bD�"�392�	���Ҋ:u���b4��5xx�����q��
�R	���~��Ԯ]�Z���S�,::�QSK_n�WɌ�����S�NJ�I��i9���ݽ�++7Ν�BKK�A��ba�\�K*�B�`�4;�<y���T�<)���IT�,�?�e\���W�Rq�z�U+���T���c�����1��3�e~��ի�ѧ�V܁���D?(����1i��1BO�����_D�#���|��סD��x�_��66#T�r|o\�Ν�Ĥ!�00����������C.W���G޼����/��q(�'�U��BW�Ϟ�B�o*�\r���XN������ޯ�ӫ�_��G���ʲy�EN������W/���d�8�o�ĠA�(V��"��'��ʛW��K{ѢEu�O?�ݻl�6��5�S���f�����,,vs���Dw4��a��}ט7�8g�L%�@����ŋ�,mٵ�
����+W4��R���z�1�v�T�B�GԨQ����L��
d���@LL~~A>|��/�����2j�jb�jE�w!�z��˖9`h��ٳ�$�<~:}�6	%:{�+V�cɒ^�PʚǏ��Ç���Z)�	����!�:u����L��415]���7S�F��9xp���L�|0���%Kz���*��Bڈ�G<z􎀀LL���Z@@�ξ��:�Sw�Ǭ[w�?��)�
YN�ʥR|�D"A*�P��6zz�)S&*#��{F���A�*�]{�ȑ64m���G�0|x��Y��-C04�e�w/�ɓ2lXs,,�+eM�\���17o$J��A\/��*W�(ǎM`̘�̚u�3���8%*U*�Νøp���k/$zLݺ�<�K�:��Ѕ�[���ٗr�R�v��^۽�*:������L�x�.]t�v%i��s$���ϣGA��I����Ls�TBɒ��;׌^�2dp&E-�GddǏ����� 6���̓15�e�(  �ݴhQC�=���=	e��QJ[S!�SW�2{vgt�4�����m���p�fUY��7�g�nݲt�����ٳ;s��=6lpfΜ���r=��H��K[�¾q��m֬鯂���{����_�T��˼~�	/�Wx{�NHp�y�	�b�
P�N9�5����-ر�2~~o]G]]J�<̘a���q�O	��������-��e��рR�~yU��ㅆ�3p�*V,ζmC�ݬ�;�\�����݀ʕK*eMA���C���??��í11Y���UK��jƃ��2� ��S�Q��!E�`֬N,^lπM��b%I�T
��޽ &Lh��k��7)R$?���*�,�֭��ݻ��O�P�|�G���'8������?F �J�Z�u��¢9uꔥN��hk���w��ɓw�����C]]�B�ȑ-�<�C����[ED������uˉ]Y�B��ʕGX[����G�2E�8�6/3��Ѵ
���{G*uį���<	f�nK��)���T�\��L�~����1o^7F�n���/]ڛǏ�6�
G�hi������[ۛ,Xp�}�Į;eI�Trs{�T*�)�+��ڍ��[����Z���=f�g�.�M�z�T������s�^ ����������2����W�
�Mv�5J'4�TW����T�y��(_>�6��^�ʏ��:��Q�nݲ��렯���^�U+�T*���ׯQ=zkk7�?�@���عs&&����@H޿GӞ<9Y)�i���l��ˣjՔ�MAȍ
����Cٶ������%k��KQ"ZCC�]��ѩ�ZƏ��޽#����KY��}�l��%ڴ����J�!��t��#5����s���9�A���(����!��G׮zj��p�lL&����5��/���޽@C�H$T�Z==�T'8S��62Y�C�J,^�+Eɺ�G�ңG�4�39
����p�χ�V|I�ׯ2
TSVR��ѣ������Eܿ���+��^bk{���X
ʇ�ny��t00�AOOG$�2�ӧﱱq���;��
z�n��ݖԪ�s?+!�-_~{{Olm�$�S,=Ν��ѣwl�n��uAَ=����_e��D��S55q�2�D"a���ԯ_��c�af�+��T�X<���,Y++Kz��̊�;���͛W�s�����iZ��!0(�Hz�����XZ���ݻ�ү_c��4UU�)
f�<��fV���p�l�ݻ/ܾ�"!�������X��O�17oD�i�@��WnbhX	33}��o��x�ʕ��d���su����[�<y*�7oe$5��J޼� �����J;gNV�Je�U+E�j��ӧ�H��{���/��|���;v\&.NNɒ�v�|�"�,�G.W��⋵�;nn��X�83ftb��&�������{�-[\ٴi��Օ��B�`�:'����^��R��Ԋ���w����W������E�vg�H��J��ϟ����#���T���B��hQ'��aM��kٲeH��M��uX��Ӧ�Q�~y�u�����s�h�f%��bРf~�!Q�N)���;Z�^�ŋ��]�l�����h�n�/��SC����Ɲ���$�NM�а������O�s��sn�~έ[�	E]]J��e14���AE+Q�r���A.W���;�_����o?��7��Qxj	�P W��J����Wxz�'C^�@G�xBD_���O���˗H��޽�x��#�Z�d���m[[��؅>�a�o��2qb;����ƌ��ŋ��Y3{��9ǘ1{����險�.E*��P(~��~W�nYΝ�.����EG�2{���˜9]?�����Y�����~
u�����Obo�k��{�tI�Tر�2۷_�޽?|��3�~~A�<9I�ѥ������i-&�c�U�#d1��r||^s��n�z���/'�<4hP�&M*Ӹq+�?���er�� �_���7w� &����hhH)U�0��ӕZw/$��ǈ�ȃ�ɐ���&�z��	�At�]���A����[���9q�uu)}�4b��T�":�g��ҧ�V��m����J__�Pо�j�W/���C��� ������_��x�TB��ظq���/d);w^a��3��ט��͓�߈��3`�vC9wn���?F`d���#[2sf��=GI�T0`;�څY�n@��"#ch�`˖�ӫ��
�K���X:w^G��y8uj��`�����}����]{���/����x�4lX��M�ҨQetu+d�f�����4X�O���MY��o��������b����~��^r��K<x���k�~�"Ou��+��^�n��T�R2��h�����荍�7n<�Fm�3�ܼ!�'IYEP�gLM�S�Fi�!����5��Y�W��R����Oѱ��~���_}����%9;�2a�~tu+�{�e�CC���e=::Ű�����֭��Y�ĵks~�f(��Hz�PT��:u�n� �w7H����M�.u��c!y�f�)����..��P����T@��/׸v�	��O�y�9_�DR�d!�5���qu�4�B�j�r\�Jr>|�����~�f�jjR���*��^H?�\�ӧ��y��g ��oh���_1!R�lU��T������d��k�F�u>ܘ�ͫ��Ƴ���(z���ɓ�i�
����P�JIv�L�33ۀ��K���I#�J<�˗���[B����С�ȓG�FQ��wP>|�3�܌E��i�K˖�12��Ãw!uD�#�\]���؍����u���hҤ
tWat���������a�@���:!�����kמr��BB�)\8?FFU12���q����f�ξXX�N�{$	˖��¢yE%(�L���Oϗ<}���F�ߛ��P�h�k����+ll�8u�>
�e��&XX4	�,J&�cР<{��)�)�1ɷ�<�.!����Ō���?�H$F�l���}��-����íx��;wZ`l\�ǟ<y���k�0LMu�~��}&L�υ3��!��Hz����w�{�qp���5o��t괖�W�6s�~��m�UV��r�o�b�~���~\��G@@
�i�*U�y�jԫW>�l�O������� E�-R��1cZ3~�L�L�H�xy�N�r�~ �^}�b����[]�
Y���L��������Hݺ�>ܘ�=ɗOC��	IP(L�d���/'ONV�h���rmۮ�N��l�:$C�!)�ƍ.;v��E���Ǐ'�ǃ�w�� du�ѱL�z�s�X�ܜ�����?�8�ɓ8:ΠR�@���k��,��Ç�eF�9�Hz�P�V+��M�3�i"��oGy��G��Wad�3c�a\\|�t�71�1�����%?._�����dqԭ[�6mjӦM-6���{r(��G l#""�e.��j�jU�={F�����ǈ�����3$$55)5j���?H|�U6Jc���8p�O�"�ܹ>��-hҤ�J�Rg�2v츌��-�;~�.Ӧ�q����n������{6mr��	ʗ/Ɣ)P(̜y����D"aڴ�����m)
V�vd�zgƌi�ܹfI�/���bf��B���Ԅ�	�o?�G�M80��mkgf�9�Hz�@P�gq�䤄ǈ�h���zu�z|de��~�+��t�\_��J����\��˗�	
�L��iժ&m�֦U��b�H�8��o��T�B�x��qjT�TG��hjf�'�B�y��SBI���K��^M޼�n��'��޹�kk7Ν�H��Ԍ�C�Dӳld˖�,[v�M�ehc��X9-[.�iӪ�]�?��#Iy��7:s�'�*�`��t�� uu)2Y.�Ç�@|����M�4������;u�Ӧ�ѪU-�m��}c``(&&k��݀�+�$|}�H�={���,�-�D�#�����G��_���n���Zu�{�f�ч_�DҦ�*�7�ΦM�T��N�_��.\��ƍ�(
6�L�ֵhٲ��D�JEG�2�	lmoR�|^����vaBB�+GMM��dMMMJѢpr��au�B��Q��竄� >>o�����ʇ�n��$���N��FE�8y�kkw|}�``����-03�'O���X[�O�N�d˒%���4��s���`Μ�\�6���f���>|ˆΜ=��5��2�ff�?ݯ��q�E�N�paF�n��p!Cxx0t�n*W.��}���y���͈6?$�_��@��+Y��7�7�̰�=��H�i�����1	_33[��a%.��wfS�����\�<�=6I�z
����p�gg_>|���&m���Ĥm��FKKS�af{o�~f�Н<{Bll5jh�xqO�U+���2�ã��P�y�j\���D�ٳS���Qu�B��Q�!O�#�+(U�P�n��=BR�(�ի���{;�[DDDcf����-00?�ّ��/#G�0fLk����~11�-�ĤK����s	�w^^�X��''��)˴i�ԩ~�g""�i��O�O7a�Ȗ�� d���?0p��ե�ڎ�b���h�i�����ө^�4 �����>��sŘ�TI�h��O,-�?�-��jl�g�ԭ[N��%���}�FѾ}U�#�PT�7��\�����/��aT�X��ұc]�4��-vew�<g��]|�C�|y�3�+�7K�r��m�M�㯿�Ү]LLֲjULL�8r!�	������1��V�T=�
	��z�ʓ?
׮=���gg_J�,�СFԌ�%��;��޽@���J�ކ�\�'�'RXY]e�RnܘG��Zz.A��dÆ��<D__��S;СC]1yE���2d�N����o�(tu+�t�L����|��������çO4k�c�ԭ[�i�L��bܸ�(�燡�?D�#!-��������0�\y''\]g�8�䅅EѺ�
Z��)f;g߾���ꇽ�.^|ȷo1���`bR�ꊱ�d�Z'֮uD���0g�Y��?��ad� (KHH���������F�%K"2RFXX$��g��6t�'��ٜ�_}�n�аVV�^���[M�.�ܼ��2%d(o�׬Xq�K��iذ2S�v�!��ьe�ݻ��5�֭k����O̜y��ןСC]6n�ׯQ��o���5 ���9�'���˗k���D��G2���%���.AMM�\��i����Ώ�l��#89�p�����Z��[..9{�..����Ȩff����Oq3Phh8l���e���z���U� ¦M.�:u�LN�b�"22&�Q��~E��*``�(U<=�>��>ӵ�*U*΁�3�	�-ٰ���7��mB�x��+W����:̞ݙ�-k�:,A��d�8f�<̩S�X��}�4�\��/��ԩS?��L�Ў�'�Fl�?�����~}n¨[���Y2�]{B�fU��ܼ����/��q�Օ���g���d���"��DF����bi޼:���sg]qC��bc�����������2d�+V����J)
��ce��ŋ)[�3ftb��&-Z �\��'�	cs=<ط�ڿ�����@G4�͢BC�<x'E�hbc32S_�F�e�+#G��A邃��f��ݢJ�R��mI�N��5UR@CC�����]��S�x��#G�d��]�������/ǖ-.���Y�w�����"����
zz�c�Ԏ�H��iVK�v��^�466#T�@|�|9}�>/>$.NN�����U�Ν맨���~ׯ?�?����{�եl�6SS]U�%�b��1;vkk7?~G�fU1�%&&��-y�����y����|�ӧ�RK����Q�?ScD\��}��O�����s���LKL�Xq���op��<���e�9�����H6o����ŋd��N��7�4!�ll�Y�܁z��q�n@�n���DGR44Ԙ3�+cƴ��H���������Q5 �f����X�'�w��ڵN��|�ر	�%W��ܺ��c��r��'߾�06�βe��ԩ�� ��޼�ĢE�qpx@Ѣ������v4TTuhB.��e({��s��-bbb��ӐmۆP�v����������[�ã��z��$�����Zu�o�����
	�R��'��1v�>C����i	���/��u��~3	A)"#c���ʖ-���K��.XX4��!��5��e.]�KHx )Jx|?���^�&~;����O(Y�5kj���@���UV�>|���X���څUN���ĉ�<y�7o>ѠAEf�6�[7J�(���r��([���y�EJ�֢N���q��x�VP	w�'X[����K��ZL�؎��*��`��UKH�C|��v��d�Fg>~�@]]J���	�b��u�YS[4IU2�B��ivܸ�C��e����r�D���<��)�L2Y�d����G3vlkƌi#�f
�(
�O?����O%+)+��?Hɑ�"��nnO02��P�x���t�˔�۴��̜y�*2dH3U����ԩ�;v_�7T�T��}ѻwC�T)���r������N��s$S�t���	��A92N$<�L��['Nx`e冿M�Ta��!t)]�K�(H��u~[���G���'r��}""�ɗO��u�%$B��*�F��l�Y��=������?~�x�1    IDATǑ#�Y�~�x
/��\��������y޼���Es�N�(���͟����"����ĳg�Q�"��I�^�0gN ~��ի������~�����������5���r��������*��=X�*�*���;��;ɵkO��ː�~3e�������ȑ�*��x����%,7����g�l�0���U?%�B�bT�P�n���fhO��O(��o���� �$BD�Ԕټ�"۶��q� ���g�W�8G�Ze�ѣA��W�9�_��x��-���5k<��UuX���\�臵��R���1��_�(TH�3��Hz$�ѣ �|��I�* �;�E�bh֬��#KZhh8˗�e̘�T�VJ���h��A������;DDDcbR++Kڴ�-���PX�7֬q��ƍZ��p��4�a�$[<=9rd<uꈄ���n�x���U��|(Y�cƴf��f/�u���ԤԬ�M͚�����O����MH�89��e�ńF���ߧ�TD_���>E��g�5�/?˲e���+s��ݹ�GGo���"����:�_b����?�M�6�pu�M�ڪKr��M�0n\����o1��r�3j�ٳ����$`."��$��ƍ5k���^�D"�w��Ԩ�����-IS��ƍ�\��{�.�ɮ""�qpx��7���J��ؔ�}�>*&�+8r�6K�:�P(��.��T�س�[�1���U�]��d�<����n����a�ʌقΝusT2���(��^���˄�ׯ?P�rI��+���#�^�r��zt���M��?�0qb�L?�n������q�~n!����f����q��勲hQOڴ���!W�������l���۷��J����� �$'�H�6n����N��H­[/hܸ
����0n�z���TV�n�|Ʊcw���ko03���+���3������T��s�ҤIQ��xx2o�q|}�0thsf��& ;v\���M%�ʅ�����	%,���t�n�ڵ��ӫ���2D�B�h޼͛��(�Ç�7J}�S��5�&��P�f�L�c�J���̘q�)S:�$�q��78:N��s����+W���7�g�2bD�����.�<XZca�''�nu��# uu鿦�(�J%�ͫNl��,�5���x�T���/��H­[�7� g�>�D��Y��E&�cΜ�o_���:�!""��G�r��||�P�vf�6�W/C1f6�c�r��K�fUqq����[��,Yb�ܹf��)���u�9VVWqt��x�ђ���Q�d!U���J�,D�u�Сn��^�M(���|����4J�W�<���!�+��1Idgg_&N<���-�=�s��?6V�����a�%z�Y�����A܌�3;�&���BR��Ν�ӹs}<=_�m�%Ν{�D"%66�BA����V�ׯ?Mh~��&E&��L!��!8�KB?{{O�t�˲5��v]!00��{G�:�l/  �={�9t���rz�h��}2�۾�k2YVVn�]�H���ٱÂ�]�~8��/���ӧO#Ǝm��@�)::�S��aeu�7VdÆAt�'�����Nqtt�ӭ��(�ɓ��� �o�`���R5�N���Ɏ#���3z���m��U���M^��ȁ�Ur~!�x��K��s��}ڴ���̓E�A�b��uرÂׯ?ac��޽׈���ݻ/ؔN��h�id�8��U'22���Uv�#zz$����̛w?�e��|�a�E;6��M��N���Ң�2&Lh����UN��P(ps{���/>�|�bXX4gР�	eB�p�?���I޼����m�8���i�pLXX�:�A[�0��D�x���߽an�33}F�h���h�11�����{l�+�����7J-��~|�T=�
Y�Q�;/��;����_? 5��/���5�-�ѽ{-���������.̢E=~إ%��̛7��K�*m=�$���EK�2Y!!�QW/FɒCQ(b�H��4�W�93�ܹsY�dI��C��H�͛�hذ��RP�d!7����l�=E�O�� 2����w|����W6BdɒaD"�,{�Ѫֈ�j�h����h��jUu+��"��#V�EDȒ=e'�~�\Q#Hr���|<<�u�}G��}���(f����Ys���$:uj�����ݻ�Zެ
O���_��ȑP��o��MS�����<�B���JX����^�իQ�^�ϡC�11��;�td̘�XXT��򠯯����#�t%�R��c�cݺs$$d���E��$BZ���O�S�]�c̘�t�欶�(��J$rf�죖��o��@��z���!$**
===|}}��~KZZ���  �)��hiAVV1��[��x�eԨQDEE��qD��	.]�˰a�ekˀ���ömW������_YZ����^B"�1x�+V��iSku�&<��j���'i����[�ҩ��S~��8q���?��ՠ�f+.��{wk֜�ڵ8��������!N*����K�嗣df*�:;[�����n���U�&n�HdԨ�xy5`ŊqjKx�Ʀ�r�)��r�FW���ļy;�p�Ç�e��bn� Tooo�����Fڽ{w�G�)?&99���4ڶmLbb�̝;@�a��\����wХ����Pw8�BHHK��Сk����G�9��L��
{������-b޼����b���|��@Z�nX��
UErr6�֝cÆde����n,\8//1�Gݞ4(5&��A�AA���@~~1�j�Ӳ��j>���vv��Wtt#F,��يիǫ5)�p�~���3���b4O^^?�|�ի�qq�a���bN� ՎHz<�ҥ��rۍ/`jj��'P۷_%<<���?Uw(����,]z�[��ٱb�8��o!ZX4Thh<���zPqՆy�<�j#/��?�@�.��n�
�T�*bX�Ɵ��C�[�&�Gw`ܸ�XZ�;4��pp0��7��R�R9I����W�#��13�� 	⠪yի���e2dȟ�ښ��ߓԺ.���������V�u�B����W_�H�=��FV.� �7��x̥Kwi��]��OW�{���)���1n\G-��F��9ʟ'00�N��زe*�;?�5BP���<�,9���pw������ٕ�_~����"�,y�ʬ�ʗD"c߾`||�	
��E[~��m�z�C�VR���4kfC�f6�����b�_����}�~��0�L��l�����ՖZ�J��HJ�ϰa�055d��)ԮmPn���(
���M�n���ᢶ8�!ZYA%��=&  �����]���\���C��_=�L���O��;�#��ع3�e�Np�N
}��r����ņM%��ٰ�K�BOO�%K�fذ֥N^�<y�͛/����WO��-%%���ϳ~�923��߿_}��FV�	��fM}ڴi��0�<UKLHH,�y���\tu�qr����OO�|��+'��s1bzz:l�<#��k=b۶�������?��!��heAx2��xHAA1���L�֓S�n���M׮���qq�����o�u�)((f�Ƌ�Xq���l�b���4ib��Єg�p�����֭$&N��̙�^�iQ��y�v0x��X�'<Spp,>>gػ7�:uj0zt{ƍ눵���C*���!=z�<R�APP̃!q��H~~15k�Ӣ��jcLÆ�|������ء������,Zt�1c:��d��X�*ie),�,� (iii�P(����]d|��*3��xHHHR�//��v]�8k�*��-\����1���C���֯?����W�ȑ�2����w���9����}��D�n�,_>�ƍ_�U��ߏ������o�C�Be'��8p bh޼>�㭷<10/¿��L��3e�@�|�LNDD�jm�s��Ys�T�����5f�Ƌ��)�c��Փ�X����Ţ��s'�9s�s�|$o�ݖy�D+� TWOKr<��#U�x��������17�É7��7��#cط/���߭�C8%�6]��_�r�~��wb���j��&<[Q��+N�t�q�իÚ5�������Ν���R�	���RSs����?��#==�~�Z�s��k�Xݡ	����6..ָ�X3bD;��s������F�hGtt*;v��OG e�������;Z��+�|������'�=�5LL�InuS\,�?����89Y�g�t�iJ�)D��!���xy9p�r99U.�P(���=t�ԤZ*�J�����?!11�1c:�ᇽĖ�J�ȑP��z��9L�֓�S����H�B��9�i�Q�ڗq�Beu�Zk֜a�� 5���u�_�+IM���{��R����[����	
�U��]����9��h��d�����vxz:��l]��U.܏�U]Ə�Tf�)Tg���϶����ܹ�0��+�A�|J�N
��.nIy�M��*4�t��|OS���Cbxｮ9r{��x��5�9v�u��r����������Ĥ���m�����d���La��]�:u�7������x��e���ŋw8|x��Y��$�]g�j�^���ņ����^מ(T>�����L�ΝӰ�������kѽ{S�wo��ڽ{��$HPP{���WD�z���1�A��ܹHv���w2zz:��;
�Gzz.�|���ۯһws�n}��_OA(���xƌYɰam��ř6m����fn<)�P(��y��_5�'����i��x 11���,����s�uw�@"��p�~�k�����éP
��c����Cܺ�ȠA^�_��K�Q*Nnn?�|�38;[�}��o�����~8Ȅ	�i֬z�{�������E���,��9������С���C������--ر�,-�>�F���	��&�(�ܾ�LH�rm�ŋw���H$2��k��a�J���?���D"c޼����d�Pu)
�l�̂��QC�����B�a	B�r�n*��٬Xq�?��C__���ӽ�]�8Ѵ�u��$��*�ܓ)����O���1��頧�Gtt={6SwH*�֝#%%�ٳ��;�
�_�$$$��_oɲecpv��5�B�`��+,Zt �D��_b̘�e6����"��yL�޻L�O�\BC����g��@j��W���ٙ�;4�
IL���{::�l��/_����MӦ�4mj��o���BC�Zcv���_��P(��5y�ā�-m14�w������2��}�OA�ݾ�̧�n���hƏ���ٯ=�x�b�����gP��9s&�s�n#��155�gO�vmJ�NN����<eQ���Tj<kˋho�D�qu�υ�����R>ٺ��_�����]K}������d�����D�NM8|x&-Zت;,���cU��ѣ���'��t�|Q���?ƤI]��jD*�s��u֬9�ŋwh�Ԛ3d�5k��H�������{�l��~������� /���ݿ�Opp܃չq�\y���|�&M,qs��qc~��(|�C�wVq����Ï�K���bÁӲ�����j�nݚ���\�@.W��gd�kW۷ и��{7##� ��2��<Ok�y�1E{K%��WN��I�n�S.�z�?��2�N��P�]^^K�篿NaeU�ի�ӿ�(߬��sY�p?[�^�m�F<8W��e~�u��QP aʔne~߂�������"��s���,��qe�֩t���Є*�޽L��CC�n�Z���֭E׮�t���ZBBAA1�ˎW�J���'O�T�Ɣ�)��z�9�g�m'55�/������>AP'�T�Jn<��d��##���L������~��:�Ϛ顩D�e����q�ہu�γt�hu�(��,_~�>聑���U�\�`������A

$|��kL��Yg��R9k֜�矏P��K����7=��w~~1K�g��U�߃ 7n$��s��;���eĈ���	{{3u�&Ta����'u��b˖�eZ���ll���1����8w.o�?Y�xzz:�r�J��s�DFݺ�pw�{�:�ww�r-��^VV>_}���[�п�okk1�Tʒ\� 33����G����GFF�����P~/==���:���62������׿��U���ᖑ'��<o�ʫ&!��x�1E{K%�@Q���")2��.]4�*�e'���a���ܜ?�W_�����ri���ٳ|��.��Ә:�;Ӧ�,�>�u��#�ə4�k�CP�LΑ#��Ys���#i�Ē����ۻ5�j��|��(���l�<E���$��^:z�rMw�|��b)ׯ����o_0����bcc���������fG��b�&ڳ'�/�؉��k�L�J��$���dErr6���瑖�Cjj����Ir<�vm��jcfV�Z��Ұ�9&&��|��[���ituu���iӈ)S�ѳg3ƌy���m'y��K�s�z_����I $$��ukq�f"��q955��P%��GG��`�^�N��MY�t4NNbHiep�^&����С������O,�m:r��u��1iR񆽊�?_���IϞ�ؼy
�;;�R}�BDE�2t�2�իÖ-S�[���C��3��f�a��������倗���k����*g��Z�Or�}���pt�|dcL�f6��R���3gǎ�1jT;>�| FF5�� ��\�P%1��sIM�!==W�'%%��=^�������!�浩W�&&��ۛbbb����2����}42�Af��6tu����f���L����7�T����D$=P&=���8u�&�{�; ~�������Aݡ�)�DƊ'�嗣�ۛ��;Y�ܫ$J��-_~[[�
�w�X��Y�۱B�'���7Y��;v�����o+[X�:j�"ݹ��С˰��˦MS5�d3)�>?�|��>�U��FF5��ř.]������Р�X�FNN!����hQ7��4jTO$˙B�`ݺ�|��~�իöm�B�%��IKS&-���KJJ6��9��吜��Jjdd�=2?CGG[��033�^=#Z����Ԑz��`n^[U�an^�\�Ǎ�j�����(r�����]5�]�U	V����D$=Pn�hӦ!��� �.��e�a�~���J]}	���O��ƬY}�<�;��b0We�_������2s���z�֧JN.Wp�h(k֜���7������ۻ���*\hh<�F��J�kb���o�R���+4��6���X5 \.Wp�Nʃ��X��bX��<�#��xxثZc����e�Muu�N
�|����h&O�άY}�QCO�a	����#5U�F���MZZ.��ʤFjj���IO�%--��DF�zXXaaa���!M�XҮ]c��13�C�zu033��T��Д$lQ�T����-�'w��Z����Ht��j��(((���$��`l\ww{u���?��ޔ!CZ�;�2��]ȢE�Y��<;6��g���[Iܺ�ļy;�p�Æ���^��ҨBc��H�ܹ�92�B�+����6n�����޽�uk�ƍ����Yc���˕+Q��
77;֬�P��^ũS7ٽ;�M����_�oٴ��h�Ē&M,��n(烄�%����|[[�� �DH˖vU���<I�r�-;�/���ɊfТ�����GH�r��rHH�"55������f���EFF))٪����m%zz:�����R�̰�4���sse����浱��[i/tL�܍#G�3�[���ҕI�Oz��' �ʹw/��]���V�����o�²ec�DġCי;wR��_�СU#�S�eg�x�!֭;G���ٻw�#��i�jZ�jP.+p���Ě5gؾ�*::�x{�f���4lXOݡ	��ɓ7�4i-]�:�b��2O&����bf��Ɛ!�*�
U__�A��=��+���]@PP�ju�'IM�AGG''+<<���T&B����jէ	�c֬�ܽ��'��ծ�Z�Te$$d���Mb�}RR�IJ�Orr6���IM�y�*���#���R�^-�����ym,,�P����թ�ո2��O>�B^^�������ӷ�UK�Z���S��k�P}ndTCC�� ��J_���c13�M``��Tw8,Yr��M�y�����$&f1w��cذ�|��@���/�5��    IDAT�\�`Ӧ�|�����X�xÆ�Q[20?��ݻY�x�Z�/�8�\��������̙40g��x{��N�l��}���6m�y��O�5������W�W_���8��jҵ��#��{�2	�!$$���Xv�$?��Z��i��N�-���[���!��
%���!V�:M�6�8~�"�+�����IJ�V%0J���Y��䐘���x�2�vm�����T&4�4��ʪ���551\��R9[�\@OO--�k�B
����]��֭3* J�Y���8$$�ƍ�q�r:4Qk,������Uڒo�\�ڵg�ᇃXX�u��t�(sU�̙���7�0�33g�U�&�Ç����%V�U�مlެla��I�kWg֯�nݚ���N 6n�����x�N|��[�:{��=V�<��?�̬����[[lmM8�P^��H"((���N���ʕ����ԫWG5 ��5Fݯ-%  ��?�Djj6�}7�Q��i��N�L99�$$d�Ibb����w/����$&*�^X(Q�����2q��逵�u������66Ƣ
��һwsN�G"��Jr(ii)�"�j�04�=���U�����ؘP��	fj��кu�J��$..�?�%((�>����10��1����ͷ��c�� :vl����4f}��Wy�u71�M�ݽ����?[�^AK��[3aBg7�Pwh���b�),�ˌ}��~��Jʨ;tp�4-�::ڸ����b�ȑ� e�޵kq�֘�/�x�!���hԨ������W��Ujp{Iu�_��kWg�l�������4PAA1��=���$!!���,�rr
U?_�Nll�U�-��5���TU�aii����ݮ
��u����R������:,Y2��[��q�F���W�A��")IY9om����L�M||m���EG��	M�m�6F�Y�ǩ�g���Eܽ������ׄ]����7ؽ�C���n��_���֔Çg��b��Hd�Zu�_~9��I-V����	RRr���`���Ex�B���?�U�Ns��M���������v[�݀!TO
�����_���7y�ݮ��V�<���ɜ8�i��
�UK�v�Ӯ]c��RSsl�Q&B~���������ZwwU2�����fƌM$'g���>�m��=�WW\,%>>����$$�$3��Jtde�~�fM}lmMlZ������u��V&9ll�E�����Bi�hkk��Z���z[[���#�H��g���#9ِ��Z�d�瓒�GN�>!!ʖ9c�"���^�X��ۛ�Ç��q��x����'���|���~���by�����h�q�d���2�����ӭ<x�����g��.z�*��'o2o����3mZO����US�\y��+Oq��=BC�}�UV�����d:uj�ĉ]�ݻ��$h�D�̙�ٻ7�_ɠA�����2���>��Ӧ�Tw8�N�Pp�n�$H,��1���Wʵ�%�+W��sg'�,y[TwTq��R���$..�{�2T��e�AJJ�j��.66&XY��������BC��drc����/�����$����(�1�ӧ�y�A�ii�����牌LAOOG5��С�4o^��>�C&S>�bb�T����T��N���111$33O��AA��9Q�<��o1}�&tt�ؼy*�:�w&��|��i|��.���0��m�ާ~}�2�c�U�'� !!��k���{���b�bŊ���K�XyyEL�����h֯�.]*f�ɫ��m4h`�����J���Ңqc7�P��K	�WI}|m����jF�����aƌ�$'g��ތ!�;��DF|������<�Ԩ]� ;;SlmMi�Ҏ�_w{�2�an�y�y�'�?�ӧoq�h'O�$33���ٳ������@X ]]����q�i�襏-��9u��ןW���d�v�D���C���N����/ܸ��L�@GG�~�Z���3T�Gxx���TOT���Gi߾�+�#�HEER.܇��tgѢ�ԭ+�Ӛ,/����cŊ�4jT���?P{K׳ܻ�����������Z�r%
���Y&O�Ƙ1��Z:��KM�a��U$$d�}��li��Je׮@��#ػwz�~㪯�������6��H���ѩS6o�;*�DFBB��R��F\\���U�[���P�1�+�۷�9v,���ùr%
�6m��=���GG圲���l���-���Rз�+?���Ki��La˖�l�t���<tu�UɎ������dI������Q(������]]T뤇��R�֓�7��g��)j��E���3m��X�tt�(��
{����{((�0�����K��ۑ#ױ�������C�v$���j�iBB�pw���F1`�[�>*���4F���={>�As5GT:YY�̟��w��$����Yks��c��6��*�<��>\ݱh�PF��Y4QNN!��iDE��NTT�ѩ��f��t_u�X��>vv��ۛѼy}��k����*�ab"��UIq���11阚ҽ�K�v�[��OL`���cl\���tuu�����0bD���#44�q�V����H��T��m/��Z���`�>�N�P@�./CuQm���[�����Rk[�o���ݎΝ��Ci(
���4��U�l��ƶEJ���̛����hF�hǜ9�W�+�_�O���dJO�e������9��sy�|��`���;4A(���X�yg566Ƭ[��F�x�_���@��>{MݡT�Z��xuǦMS��!5��.x��H#**���4��U&7�Ҕ�ut��_߄�qr��g�fUj�j�jh�l�����Lr��G��W���zлw3<<�[%���E�����L�&�\��+m�ۿ?���,����<LGG�"**�?	 W�����9�m�#""	�T�T
�۫���Ν��a�ډj9~ieg��Ǜ����O_���{�9,##�ŋ�a�<<�9|x����V�ee�s�r�_���i���V��g׮ j�2`Ԩv��	kkQ�-T{�1c�&:tp䯿�ahh��J�ȑPv�`Ӧɕ*nMS�������6700�36��t��ʨQ����dd䩪4��҈�IW}���(ׄ�ښҰ�9-[���n4lX��ͱ�7ՊՌB� $$�������ڵ{�ұ�#_|1��=]^*a9sf_<<�8��+?�f�~�����F*}��Y�L��Oly��ա_?�پ���m�#44}},,����t�q����ի�Z�_aa�L����b)۶}@۶�c�Hu$��ٰ���fM=~�m$�{U�7d~~�%�|��
�e�jΟ���ي3d�5k�(� ��B�����oǘ4�_~9���9����<f��ʘ1�+Ͱ���IksSRrTCR^������k}�����6��ꎎ���;�\Zf����\��STi�[��Fvv�Ll�ۛѰ�9��<��Ӡ�9���߾+����"N�����78~<�������ի3g��S�&��>���
gg�2�WKK��~ITTaa�Olk-@��
P��h򹤦��I���xj�ҧu�j9~\\;v\e���{R�q�E���A�VX�ll�*�nΟ��/v�̻�veƌ>����ѣ�t��"V����B6m��ڵg��l���S���Ic���i��>}#G�����TW�+��swP��>_|1PݡTu�ݻ�j�ߓ��n�p^�6�q�z��fPPP�ܹ�2��x�|r����"#S�};���d""��};�����@tiذ�ӡ�##G�����̩_ߤR%6������8>�L���=��w�g�f_�����cy��IO�}B5Ǔ�%LMkk��	��YEX�=
��j���ǲe'pp0g� w��Y�R9������2}zof��+^`4T||&�c�� �wo����J3��I����<y�ŋ��;�*%**�5kβe�% ���0qbg5������$&f1n�j�زe�#W�+���Cػ7�m�ޯ�I��iks��b��#�9s�5�(,��`�^֮=��������i��\M#�ȸsG�ظ{7�[����L&22��B	 VVui��WW���тF��am]W$����J�\�|�'np�h(��)ՠkצ�������R�f�ܽ����>� 7���B�jk���65j�R\,}b����}���/�Pm�ׯ�SX(QK�Fr�}6o�ĢE�7#++�ɓ�!  �+��������P�_��ߎaeU�u�ޭ�m��K��SL�~U
���go�z�?Ǐ�ckkʬY�1�FF5�� ����h&N\���!����L�!����\������4z}xu����HH�dѢ��ݞ���G��._~B#��[nn��Z#22�;wR�u+���t�R9::��ٙ��dE�.�L��''+-�k�Pj��y�<y��G�8}����ӨQ=z�n�w��m�F�rf�ɓ7�:u��v�D��;v��Sdcc̞=2k�N�����TF�ޕ��E��I���trs�04�/����|�I,,�2�U��Yn�Nfܸ�Kٽ�#Q*����7��!--�3�0eJ�J�D�$G��Ү]㗞�/(b;v\���7o&Ҿ}cV�O�>ͫ͛p�jR(�Z����֭)�9�ڵ+g�Ĝ9۩]�s�Pw(�C���,Yr�+NҾ�#6�����*ks=<�+����������DF��	���.��8:Z2h�M�(?vt���K�q#?�0���	�A[[��m3cF��i^�+�AY����x�-O�,y]���`� ��ۉL&g��!XY��ݚ��{df�Z��:::�TST�g��������|�j�����ǆ�⋁5l�ܹH&N\���>>�������������7=�?�M,-��V���;�G�Vw(�RR�}֮=���rs�4ȓ�%��B����ٳ�[�*k9�=A:t��;���ϴiHH���o�0fL��>�_�+�ʹ}��ks-,����Ã�{�L�I$2"#S�',,���""�IN���Q-qr��sg'-pr����T$օWRT$���۪����ebn^��=���{]��ř:u*uPQ���37�wo0s�`���|�����e��p�^����g�mcȐ֌ݞɓ�&::�TN۶�D{d)Uˤǭ[���jӶm�� �\y�:uj2|x�
?����q��37ӿK~�}���k���~��(>>gpv�b׮i�iS���ǒ��C߾���R	�aժ�:t�ZL�؅1c:�}�B�ϤIk)*��[�RRr�3g;�۵J>�WF2��e�N�d�aZ�j����bgg�R����쵹��1���9-:���NNV�����L�Tt[������%Oxx��	ܼ��D"COO��M�qqQnl�Ē�M����[a�	U_bb~~�!�g�ަ�PB��6x{��W�渹�i�(�W���ń	k��Ng��w�֭���/��I���_���)_~9]��_����>���]E�_�U˳�k��!��*�Gvv�}��3�b`����v�ŋ1ujw��Pi��UEr���[/�h��R9f���U���a�_�E�J_\$��z�?��1�li�O?��7=�L��  *#wҪUV�W���=���[17���ٯ�;�և�>�ȵkq|���L�ܭ�_c��67)�>AA�D�޽A��chh���%!�XZ�z�A�P�Nhh<7n$�%�)���4kV��yｮ���Ф��x=ʜ\� ((VU�O͚�t���7߼EϞͪlb���(&MZKݺ�8x�c6|�0�ŋq�f"��R�;���wC�8�3���o���hƙw�v���Zxx�W�q}}/0j�����dr��ہ��E.�;�tTwH�Cb�?׮�1zt{>���*?����0pSw-##_��]{�����oɗ_W��*''��9s��{w ӧ�f��ʿEl˖�����{�GԨ���p�=_�|���8th&..�vl+����߂��[ ��d�n%C``~~a,_~�\����H<<�i�Җ�5�����MHH�
^�����֢As\]�3n\G�6��յ~�=�4Cvv!�O����p��Azz.vv���Ռ9sС���\./�֝��/wѵ�3K��.U�Ι3,_~������߸��&<]�~�=Aq����,��7��(�TΚ5g=���{�$}�ˑ#��Y3A��^P���l~�� [�^�]��92u�Uӈ�H�o�Q�E#ݸ����?;v\�F}F�j���DU�P%]�Ŵi(,���;�����Utt���i�z����p����>�dǏ�3uj���~jo���ѦY3�5�a����2�K@���btu�i��/�xx8��l��ْ$GBBZZZ4jT{>��?nn�4kf�܄� ���wS9vLY�q��]�r�Z5`ʔn��ٌ�M+.ɨNEER���Ζ-�����̚կT�d��9|���xÝ#���*�vI�;wR����Wl���!��d��]+���+((f���t�.6�'V�i�D���~��(u��`ٲ1��*̑#�X[�����?ΪU��=���_=��C[��B�$�����#��=z���Oë�l���lgg+f���p��C����[144`�N͞�U�N:ur�S�73DE��o_0g��f��k�[w�������ٙСC��iF�.�U�BT���K�����ѣaDG�al\�nݚ��#�޽)�Ƶ�f�JH�bҤ�ܽ���O,�Ef�B����QC�~V�QV�.�q�FZZХK�^9Z��8o���m�م���j""�غ�}�~c``@qq��è0ZZzԫ7���[��^��7�������ct����P��s3e���"�l����bb��޽)������Y��UVtt|���7������ۡ�<������=�����&99�|��.�l����m��A�9�q���\�|��W�	����x���ԩS77;Z�h��im�R)���Ű}��o�B��xx���逇�����^�"T-ii�?�B�����B���x���Ռ֭V��ėu��m�N]��Ym�I�Fϟ�QbŊS�9��]bdT���h�j��w��
������#	���GT�1��]�ȑ+HH�b׮i��Rm��Fqq1o��#G�Tw(F&S�����n�q�Fv��]NU���.]��̙���Z��e�v�6n��T*gذ�L��E�l
U������M��><S�_�^Ĺs�,[v�_~A����Z�x�ӧo�����k'j솰���/G�իQ�Ĥ������m�4d̘�xx�Ӹ��SK䳲�	�!(H9䧟�������.���UCR=<��cRx!
�������/���8��th�ޑ�>{�^����棪dŊS|��>��k�/��x��!!q,Zt�O?폧�h�,K�.����6NNVv�U�Nӡ���J�sr
=z%���ٹsZ�y�������[�ah4�DR�^�ܼ6��in�qy�r%�����XZ�ᇽ=�=u�V�2P��IN�f��m������=����W�J���|>�pz���Z��T;��R/>Ċ'�ի9K���Q�R��E�p�JI�#���Bj�6��Á!CZѦMC<=�PU��q-z�p�G@y���J�\�źu�Hd��������D����,<�������9~<����XZ֥gO>��7�;;�������-��9�3uj��X��-b��u�kט���Q��VO�.�����1��Sn�Ʊca�Y3�B�����"ƌYŽ{�*�!T����k-�U	d��ٕ+O����9���[V��>Ax��;���ԭ[���?xd�gU1k�f��tX�h��C�vn�H`ڴ��e�x�0F�T� ���,U����w�q#�LN��&�nݐ9sЦMC�������d�i�F�:� ��BC�K``�6]���������*��Հ�M���=sNN!�Oߢ_��>\xqqq��������H$2Z��c������W��U����DE�2i�Z���ٸq2�;;=�F���m�������o9�VI���"��
�ԩ�w�ZuGGK�lH)((f̘U�Ĥ�c�Hx�'%%���0cF��φX��j�����jy�-    IDAT����B���0{�V��w:1oހ*y�pÆ=�Ν��0�
$�+X��$���ݞc������Zb��N�ҥ�\�Ʌw���@WW����Ӿ�#~؋֭�e]l�z�jՐV������Cpp�jm������-�fM}Z��}0�������q��Ï�K���dɒ%o?r|A}d29W�F��9n�L��Ѐnݚ���C�ѣu���:|�:�s�����o�۶�
�v�a�{�ﺜT��Gxx
t�ؤB����ǦM�X�`P�g�JwcǴ�#���k��U�֖;wRX��4۶]EOO�����/��(������W������������ukqRWQbcә>}#��1|�i�L�^����)\�ɥKw9>�������逷wkڵk�����&�,,�Ч�+}�(g���
""�V��=}:�U�����XZ�UI��t�eK�R��DF����ܤ��0|x[���j��Cde�s��M���ɛde�Ӡ�9�z5㫯ޤ}{GQy������j�?�F�c��������;)̝���S�ӽ{�r�T�j��8s&���]*�x�֝�V-}�iU!�+QPP�;��p�V;v|����(h�m�.3th�*�ڢP(8s&�U�Ns��M�����慆Z	U�T*e�޽�d2u�R�����/�N��8Ё{�ٶ-���]�v��i��1(YO�W��|�q�
9fu~\����a��pLL�1��v��Q.�j׮���r�V/*�8.]�Kjj�j�ӪUCƎ�@���xx�Wڍ)��Z4mjMӦ��P�L��ĩ��������?��g��%F9�I����_��\ `��+<x���~o�VO�@x���ݻW޿n�dkkK���U�GD$=h[	�ʕ(���m�F|�a/z�n.�^@R�}&O����x~�}�K��K�:u��̞�ZG)<�r>����h���+��A"���?�;�#5j���JI�0a��	l��~�lU��_,%���u�F"AA��������");v\e�jn�L�cGG֮�@�^͟:m_����ϐ!C��Z�ꚢ�]��[�u�������Y�fM�Vƾ�v��;�I�%s��㪄��.���DG(-�#���>���df�Q�Nڴi����h۶nn�UzV���:8ҡÿm�		YZb�	
�e׮@

��]� 77�GZb��r�?�DFvv3fl����������:t��߭*������P����pbc�13�M��My睎t��"׾�ӧo1m�LLjq���4mj�����W���M���Ҽ�U��ǝ;)��UL	��݁df�3n\�
9(_<&L����{l���+�#�l���D���ٲ�^^�Lb.%%��9˺u���)d� O�.M�f6�M�����Hʾ�Q�FQTT��0�i��V��g��1��Q<�*ΨQ��}[�ԩ�i߾1͚�T�J�acc���1� �ʹu+�� 嶘Ç����144x�{��σ�b���G�N�Ό}�Y��6 ___F�Yq�T�q�F�M�Ĉ+h�̆7���O�渻�W���˒����Q~��z���^�r�������5Nm����j��HM͡y��_�P(X��4�ޭ��4*��sƌMD�}�4q�%h4�DƎ̙�Cye���Zu�={�02���q;��D%�ȝ;)̚��	:3p�����Q�&9��^Wu���J��6o^��c�U�م̛��}��).~r�T�����'پ�*?�ୖ% UIN�EBC׿��Y�_��L����`� Ə��J��άY�7�#o��^FQ
�Rm���
%�ha[��:{�6��	����r?V��?��}���N�յ�;������
��W�����2���<�vO��������#GB)((��'r��c��X��4��G��b���a��V/5�J�ʫ���I����l͗_Tw8��q��jp�N�S��䤤d3n�jz�n��N�\<����4��(W�F��{����Þ=���j��$S����Ό��z�����ڼ;��W1���-�}�WX��?����?O����ԩb6�h��%��y����i���,���>��:ɠA^����Irs�ز�>>g��M�G�l��R��A��������q�dѓ-O ��	�/��+�)/.XXL(����r˖�`��t�֔�~����+����};�Çg�e���M�?�n��wP||&ǎ��l��r=N��GC���̙�:�{U�1+����x��)�����._�K``,?�4\ݡ�ڽ{��Y��ƍ�J�x{�fҤ.4n,&�Bu��?�س'_����WT�I���H������AKK�D�z����������88�ckk��u]ƍ��VS�Bu����G�r�B$s����]��}��J؟?�%�CV�j���v������~t_ߋ��ס_��z����N]���ݘ6�g����.�M�|�I��i^)�^�ŪU�<xKK#>���F��ظb"Buj{�lBB����]̜ٗ.]���+)m�� �������	�����;;S��7���;;S,,����lԨ�
���Ŀ�����[L��K͚���;���YJ��g2}�F�o+.T�A�Izܽ���y��Hdl�x��c;��ʲ��4ƍ[M��-�7o@���/Z��ıca��9Mݡ<�D"���V�<Mpp,�,]:��^k)Jׅ
'��4Sffﾻ�Ν�������=~��m�����]�����[���AcI$2/>���'x�w/F�:e��W*�3u�z,-����Aer��6I���<ڵkX��8x�����վ\�����С��b�/�����egz�G��ʕ���M�F��?��������5gIMͦ��|��[�jU��� T.r��i�6����ҥ���� ��M�.2�nLLj1xp+�z�OO{��G����|��z�����a�ѮL���ϡC3Y�,T�j��HJ��T*�յlʓ�f�ڳ��ߢ\��3f�*�֭���ĕ����Ib<m������W�_���Me۶+���8u��;wRX�ڟmۮ���èQ�?�3��&�M�8�ċ<�ꆩ���I��*�5�/��ܹH����R��=���Ꮯ������1X�-kO����~�c
嫨H
@ff>�֝���c��[��[�8;�M�kY<��ދ>Ο7��Yϓ�yN����!|��ll�9|x&M�X����<y�e�N��OoW��Z$=�^��M��b{�F�/�eǎ�+�W(|��&22�8p�c��ʦ�*xZ��^$^��i�-�ן�yU���pu�O߾���B�ٳ�Y��'N������s0lX�J�QF�>^6yP�Js;੷�*��������Ҳe�^H)/�:��mhO��i^�1X��=)��\(zz:H$2�Pӄ�,�-;�o���ђaÔ	�W��𪏧'}\Z?��{���ߓ~Vxu���������;�_=�̷�$'�g�t_�b��ez��?{�����w�EDTQ�`A콀�K���ލ5��h��&&1�bAcłb�{Æ(@� H���A$&A���2����r�9˝;3�7g�)�G`� j�,��:6l8G��4mZYmu���q��˞=�E�x�(`/�p��|}'hԣ%-Mƞ=W��:���4o^���Ѿ�s��mF�2Se'�����Ç�7n�z5`� �nc�u� �ʶSXۡ��N 		���;̢Eqq��W��t�撧2UݞT鍛]�Eya��	

c��?��x�ڵC�ҥ�������%����^*/_�;���q�^8�����㮞���޽����nj)2R�.Yr�_~釫kE��ST�n0Sנ���6�	�R�����ҥ��byDG'��}o��$&���Y��~돳sy��#(����ceU#��F��g�u®���rJl�[�]G�������h��Rm"�:4�&<�`�(o��Py�8��,�R�L�!�ܺ���7_0g�nʖ�T��W�ݞ
����(JV�:��Ň�_߁͛G�m;��?���g<8ss�E�i�������ڢE��u�z�j���<�`-�ٚ޽E�ru�I���g�5��g��A^���]{�ݻ�R��1�7g���)��LN�&))���յ"͛W�a�J4jT	S�֝W�|UysE�R9�G{�P(Y�nh���Um"7�k������nO��٦��|�ĉ[�v-��3;3zt[�y��;���~�g��Oպ�@�st^�P*���$�<(���o�x�޽�Eŋ�Ofذ���VT�'�@�SY�� C������@�T*��9�իOq��C�Y��'�z5��İ@l�6�G^�~�w|y 	8:ZѲ�:Ҹ�#�ʩn+��&�y-'?���9svs��K|}'R�t1M��UD[�й�<�WOк�܅��`ɒ�<.�H���C.WP����[���c`�Bevh�=�~���k�U���M�r�:4E�����o;v3]��aРfj�G�;t^�x�2�T���zD���		���k��˖��.��Wy���y��!�ə:�C�u���ػ�:k֜���Z�������j��@�J�ӓ`eU���D ��(�͋�ٴ�
��2e,h޼
�9��-�u{KA_�K�[w�m�Y�n(5j�j�������(���ݹ��n���}�E�-�nZ�r�2}�������ȪfW�@���'3s��bĈV̞�U��J�G&S0z�&J�0c����V� ������+ \\�e}Æs4mZY-)����ϭ[�ٿ��]�Us���od���(�����_'�i�y6n<G\\2�|"�u�O�r%2E���.��TT���d��� ��N�U=�
l�]�Ѽԗ��
�N=`޼}|�Ug<<4�uJ�dw��uosږ>VǇl�M9��>#�:ԑ�VU��c�����S�Ԃ�̙�L��==	۷��eK'�����}�%N� ��=��y�Q"**��ǃ���*/{ǎˬ[w����΂BGBB*Ӧ�W��oﬖ:BB�X��4�v]��؀���2bDKllJ��>A�&))���8��㉈�$9vS~����c�3R�2?�b�hoz��ϸqn�6G (��[]/YҌ�=��銫�������4��~�Y�u���Žպ���c��r�I�-�G������q�f�衎x;w^��N�ꨴ���#�={7ӦuT�ca���������Oj�))�$$�����sL��[v|||4mB�̛�B�d�|O��}��c֬9E@�=��K���]�۷1ffF�X Ȃ�4��q���!<<���8""��˗BGBBJ����FX[��@/s�2+����Ԯ]��S;u�~Q����>�
�+w\\���jղ,]�W��
��
4O�~M�ZՆ�-�
�vm�ֵ��ן1u�v^��g�����Y�@�}�<���ү_c��I'��=BB��ӓP�bi���T*ٺ��z5Pi$���4F��H�ƎL��^e�j;��2�?ͳg�<{��ۗDD���5RS�Q*�d$@�`z��M�*U4m�?����l��ʔu�T���7X��4wqcG֮J���y[�H�r"#�32�4��3Č����11o3�722�\9KlmKP�|Ij�,���%��YR�BIlm-��4cŊ��Y�{'v4i����4k��n�zK-�Q�'��n��H�rF��F*��q��"��%��{,�ŊӦMuM��o����s�>��d,Yr�իOѼyU�lI���IE�o��e�鍝]),�Y u
r�΋���XX��|�r��BCc���&*-���v�������u��/%%�=�Mrrz�``h��D��&����@��&Q���ƠmDD�3y�V��m��{�|�������X��,11�t�R��M�z�*�VPؑ�DG'���k���d
�Č�/㉎N@���o����\���/oI˖N�bFٲ%([�2��˖-�L�O/CC}d2�L�Ԟڵ+��;ԇR�dʔm\��?��"S�@ �]eʔmDF&�㏽���&�5w�/���92Md	�btZ�O&5UJ�*eT^��-�_�A��6�n����u||��ɖT*���Y�>+�)YҌ�{'�C�J���ҥ��p��*�ٳX֮=������1`@S�m�҈��G*�ǋ������8^�|MTT2��ȨbmmA�
���Z���@������T�`�����<�ʖ-�)��T*��te�w��9��h�A��n�q����"�Fj��ŋ�v�iZ�����cT�&>'��{�M�.�f�`��R��=�>�T��͛d��?����}�ߏ��o�2}z'�4���r�S�N��o��|q�zXX�o�D�⫥,X�����:45��5�^}ʪU�8r���Y2sfg>��1ŋ���GP�y'j�1މϟg���|�),��agW
{��8;����[[Kʗ��\����X�V���f�i���m|�%P�W��?N�|yڶ-�.��@��\��)S���O?}F߾�
܆��H�O��_��K��^� w��H�Q��J�ݳ�zt�梒��3�x�_��ďٚիO#��~�}}=�͍��/TT-e��Kxy�a��A�^�V(�9r�U�Nq��S�ճg��At�T���L�!j����坑3Q�ή5k������ή��y�U�X���Ѱa%��M�;�������3�k��uc``Exx�N	�))�,Zt����Ҷmuv������t��b#5k�gΜn^� ���	����J�ݺ5�O>q��\5��g��!11��~�_�2ZX�2lXsV�<������&&��1F�k)��?f֬]L��A��9SR�ٹ�
�W����X�ݝٻw�;��Z�*����)h�x�W�� �g<�&&��ۗ�ήd�5rBǎ�5m� ��9�)S�1n\;Ǝm�is�$**���tLM�06�ۛ���D����/ބ��f�r�������B�=����M�N\\2˖��wo�eI�1c'��oٺu�x]H�i�#((P�࠺�-�n� ((�ŋ{���m����aeU�&��!!!�_~9����066D&K��q�D���۶��N;Y)Ȏ��F���S��L��!G��ļe��sl�x���4z�nȨQ_P�����m��LQ㝰�Q�z����פB�RT�P;�RX[�,@�.cf���H׃T���C�����ן1t�z�usa֬.*-[U$$�����Gϳ��Lٲ�3?��eӋ�ވL�R��)^����DE�E��p�f]D��P�q���O���5mF�C"1��ɻ;ľ}7X�ܟҥ�Ѷmu��kҦM,,��pBB
`˖������냍����ټ������ϑ:�E��H�:�?�E�x�$�Ǐ�9�����+�\yJ@��|�Iǎ?3iR{&NtW�u��TΆ���� |�e'SX��p���D"��@�-[FѢEUM�+� �|��o�)c���XLM��BCcX��>>W077fȐҢȉ}�FJJ:����ߥ����˗�3��f
���P��5r�L&c�����E�%QU4i�;;�ࡡ1t��+������+uU��$99=O�.Y�#����&$�s�J4��QDF�d���_�9O��P�q.^��˗�z/�8*T�iӦ��=z���=���q��S$h�ؑv�jҾ��V�޽�*���G"�y�<��tը=w[�_?ލ/��Q[�C�EG����*)/%%��̘щ��[�,�TN�n�bjjȮ]�
��Yn9|����W��0lXK&Nt����t4�G||
�==	6WI�S��IHH�G��P*�h������ۗfԨ6����"�@u�ļ�K�x'l������3ϳ�)��Ci*V,MŊV88Xao_{{!jt���x<=�cm]<G���Y�� �V��`f���ӓ�T����:�C��IIi<x�;.s�R���r%J�==	�M^�A!%>>�S�p�x'O> >>+��k��^��M�hT~�$����Ņ�،Y��`aa�1{ ��C����/�֭��̻�����[^�N"5UJŊ�����w��4�J����Q�<�" `F�xh�]{�����ʕ�|�I=������ffFL���w��C�T�r�`!xh)IIi���������Up�իөS�"��������<��7��LJʌ��>    IDAT�:fh���])��U�<]�����4���qp���:OBB*���� o�Z/x t�Z����?z���>��F�\9�v�j�.�\�ٳ�ع�
���Kh��T*���N�<`@S!x�KK3<=]��tE.Wp�j(��������͍iӦ:nn5h׮&e���GZ����g�� �V���o2���H�١T*�4i+ii2��c`�xw�5tV�����b�u�%:w�Cɒ��*�ڵP~�=��K�bgWJE�i'aaq,\x�}�nдie��D���<w���l��ر���U�~�FRR�0`ϞŰ{�xlm-�s\'U11oy�$��Oc	�7BB�	�!%%���xq��X�4m����s#�k�ֶ��E���tZ��`�m(J��Ұ�.Ntt��30Уzu[6l����r�~8;w^���*�_'a`��L�γ�o�`�D���1_}�9�u�D__�ƍi�ؑ9s����뿶�1k�.�R9u����V��j��v��#��jQQ	̙ӕ�C[jM����8q�~����+���D"��Q5)NCCc�|�	۷��W9IIiL��g��.(�)ݰ����xy�S��3��r����P�[RR�8p-�G�k׸���IUG||r�����Ɠ'�$&f�v611�R%k�qs�A�JV8:����ZlC� %%C�	�b��q�l�	�\A`��������J�f�r�ǧ ���qn�{���2o�'FF�����q�)S�������o���(�?���������+�С-:�))�9��{���E�.=��M	��jо�3-[:�;nbTT"�}��޽��ܹ�v�ժ>���,Yr��s?�Q#��WX�Y�#$$
}}	*�~�#+||�`kkI�N�*g�\_���X���J��6�J%;w^a�?�J%�|ӝ��iu�8��ILLeذu<|���;�R�ZY �9[���N�K�R9��1G�����^�N2���ۗ�r�24mZ��?o�)n�ږ(r�����&cذ�ܿ��]cqr*�i���\��������w��N�F[jN�n.$'�ө������@=�.훯m���g���@�����C��A�ajjD���СJ����p���?���14ԧi�*�o_ww�\y��d
6o���Ň(Q�o��o��o�{^�x�ر���teĈ��sh�d:j�7~~7ٰa8:��WYJ��f�ҥK]���[��9v�.C��gӦ/ps��~[m���0f��ŭ[�4�93ft�A:@dd�����$�nE��\���+N��$��fÛ7�<~Mp�+BB�y�8���H�?�E&S �d��+gxiT�lM�J�88XagWJlE�T*gذu\���qԮ]A�&e"�)�p!�nq��bc���\�.]�Э��<������������/oɆé^�6߶\���=�#���ЬP__��'gje��@P��ļ%  #̙3ILL�Z����eCmذ��1'O>�����i4#G�a�T��C������\���$��O�;t���ѣH ��O�|�)Ϟ�һw�<�����;8���			),^|�͛���R�Ç���\^�f	T��'���
cc|}'r�^3f�p��S4�Ě5C�رv�N�P(	����(?����������=�&&�T�\�ʕ�У�+U����X�*Uʈ����J��͕+Oٺu�VR�����:�⒨]�#G��[7>�%�GWV�8�D"�C�Z��K?�͍Ub��kE~��3&Lؒ�q=ƌi'�@���U1��mD߾��J�����C�n�b�	,-�hӦ:��;Ӷmu,-��a�\_��S��l�8<�~O�̞����_s��T!x� :+z�x���^�f׮�ԪU>ӥ?/̘����M���O�m�6�w�u���E�P�dI_��i(��u�7�3h�Z��Kѣ�+����ɓhڷw��wB���(�+x�,����y�(��_��I�G��*2& NNeqt��ãU��P��5*�*�@P�H�r��b#.�e�(\]��]P��=�?��=z���d�ֵc�ضt���,s�D��s?a���*����33#RS�(�{��I��*����U^�@ ��i�-��7ϓ'O�9~<���{L���BI�2ŉ�L����]��ѬYM��A6n<Ϯ]W����L�͡��[��qq�##BC�䫬�4u�~˴i�⋼M2v��������@����G[�㫯|8y�4e��b+��c�e���;�R�y�B||2�~ڀѣ�h�~xU�T*y��5�����W<x��G�x�(��tzz��K��T�*U2�5�V��J�2�(a�i��"Oz�����s��S6oIÆ�4bÙ3�8p�&G�������]�ԥ[7���&�+X�����O��Mx�"���C��t���xx�o��@ (z�d
������G�J�蓔���])��3�4kVcc�Y��z�)�~��&�g���6G�"������/_P�l�|�u��]������[஘��̝����-uB�P(�x{�cѢ��ؔ`Ϟ�En�_��J�|��vv�����	،/�h��M��'m#<<�G�^q�~D�����+��3ҿV�P'���jU�/�hM�jeqr*+��ZJj��a��s�z([��.P��t�N=���[;Dbb*���L�ܞ.]�,��*��Ofܸ͜?���K�Я_R��q)/^�!�@�VՄ�!r��q;�o���+f�����ٰ���F�j儻{M��j���-�DE%2r�7m�Tg���!P=:����w�ѣ7ѼyUv�����B�P�y��<]?z�&n�~����|�t�4���L���[��3n��&��*eV�?Νf��M�ƾ�D	3Əwc��f/n�i��M||2����AD��a��������NNe�^ݖj��R��-NN6:����BJJ:C���Ν�l�>�:u��^gZ���'�s��-�"))WW�u�K�.uUWL]ܻ����J�xy���>�Xhh͚- 0���L�̓|��~N�|@�N��������F0�s�IM���\���qww�n]��,����gQQ�><1�%t�5"������CL�[N�z�o�����ǎ����&;v�.Ԃ�R�dݺ�,\�G͚�8rd*5j�ӴYq��c,�����0sfƌi[(�+J�?����0��¸w/�{��	��dIsj԰�ٹ�~� ''�W���RlK
311o2ċg�bٹs,�j�/�vj��'2�� ���iذ3ft�s�:��j���={�1}�N�ճg����.��4�V�81���D!x��O?e��ԬY.Gq;lm-8�6#-Mƹs�����s�eˎaeU,3L�V�Ժ�����s�%L�����Gxx���|�����<��MHHe��]|�YcZ�pʗ�$<<�ɓ�)��H�Y�Q(�:t�?��֭��fͪ�~��B�%-MFPP��q�n��Gp�~8IIi�����hM���g��Ԩa�Q�I�@��>���5 ��?�J��U^GJJ:��R7vd֬.t�\��l���̟�/�3�Ն9s�}pL�H���t��@�	�aٲc��s�ʕ˰r� �t��kcc��jdf��?� ���1z�&��$4n\w��xx8�4�˞=���:êU�U�\�}���T�ȷ[����vu�������0wn�|٠I����ٻ�����oR��
�KZ���;/�r�I�?���̘b�LX��/ݻ�hڼ��*%((�۷_p����yɣG���/nB��U�}�6��9#ӒH/&�>W�<eȐuT�d�����x,���t���8p��IO�Ѵie���;�:աL��*�� ��Jd�hon�~�ʕ���z�6I b^�x�/����2���������tU�v�5l�QÖ	܉�K���;Ĳeǘ7�GGkڷw�ͭ&�;��C�޽p�O�ɨQm�z.,�:)z�|��LN�ry����֭yJ1{�\0۶�n��B�j�>���̜�Á�6�%s�t�9���x{�gݺ3$$�R��-zz\\���ϵj�yJJ:��s��˿D��g�ԩS�6m�3a�;u�T���J�I� {�\cڴ�m[�+�d�z�6-S�8q�>R��fͪ0o�'t�T++Չ*Ʌ�;v��&��M[TA�		�bŊ���u�r�,Y��3z���VO�%��ٳ>={�G&Sp��N��ϱcwY��&�n]7�����ȱ ��M2#Fl��Ŏ���6��G'�֮���o9sfU���S�d��k~�����t�ݗP�NV����5ɩS�2e;���-�G˖�wk� ^��c���l�r}<<��~�9�^�3sfg�oU`��B�P���ϸy�9׮���A�?�:u�2V�XZA'-M�7��a˖K�׎�3;�����vbb*Ǐg'O�G.WмyU�v�K�Nu(U�\��,J��+N�x�!<<j�lY?�Y 䉫W��b�I��K�J֌ۖ^�j<\hh�P/\x�\��^={��3�@>�I�P2h�Z�ߏ�رi*�h:'zH�r��T*y�xq��*�J�6]H��.̞�5W�.X�Ƕm��>�U�ZJII������}�O>�ǢE�R���XX	

cժS��w�2e,4�ϟǰ}{ �[W��{k$8]l�[�_ƍ��:��������k�Q��=���[�N�{5�n��i4#Gzϯ�~��{�<����±cBǩSP*��h�!tt�X��%��񎄄&M�J@�=���;_|�J��� W(�J���b�	�P�~EƌiGǎ�5�h�!���8}�!�	"**[[K��3���hQ5s��ҥGX��_߉ԫg���������R��X1�<gL�q�9ϟ���隫��ߏ`͚S,^ܻP	ׯ?c��-�~��ʕ��]��-��;��+Nr��C�W/�O?}�T*gɒ���
�/@��k�y%=]Ɲ;/3E�7���Y,��J��pu��̙]�W�g��_)�͞=ט5kNN6;6���s���͛d������9��RI�VN,^ܛ�k��ƈHK���3�ƍ5m�@ (D�����{�իO��[��}���1�;סs�:(�Jn�z����166�y�*�ږd˖�,Y�'ׂ�͛w6s�B��yz>�G��T�j���_婌o�����su�R��G��Q(���7�P����
~�͟eˎҼyU�-�'�[B�r�bŊ�ܾ���ͫ0fL;,,L��;_n�z��M�>��ZW/�>����q�nR�KK3\]+R�^ſ~ڋ�� �DF&��W>;�ȑ��=�k�'����=��>���GH$Z��F�.u�رV����1�m���ٻi���+am]��
���y,���ٺ5���tz�peԨ6:��$**� |}�s��c@I��pw�I��5�W�b��J~��*ΜyH���Y3�ʕ�JAP�蜧GDD<zz*V̛k�B����6��u;w^���P��V(���Dƍ��ի�|�]�i^(��MJJ:۷_f͚S�|G��u���^X[g����w��M+s����g�+		�\������ן����>�j��^���W׊jI)�>>W��[_,-M��K�fU>zM\\�����[�?����֭���ϟѾ}-,,t3�Ej��Y�v�s�&Lpc��N��u"�J��ӧ�a�9�acS�1c�ҿ��sQ�Lq:t���?�Y�ʌ�Ɖ�ؿ�˗�S��9m�֠}���iS=KQ\�Pr��s ���pw_�?|J�~M
��r�Ήaaq�9�ܥK!DF��U*���$,�cذ�Ԭ���Ϝy�ĉ[077����8;���X�^^�NbÆsl�p���4>��1�F���?�`Æs�-[/��t�T[%u>{�իO�r�)�/?�ѣW(J��K��Z�)S<pu�H��02ҹnE 0aaq|��'O>`�Ж̚�%�-���o3���10ЧM����KF�]���q�G{����<�:E���d||���}�'O�i޼
�W�C��j�Ģ)�R9Æ���� /��XZ�Ѯ]u,�Ipp$Ǐp�����Q#Gڵ���G���7o>'>> �L�L&��/wp��~���Nz�
:�v��D��m��ݠv�
�rUZ�� ���|�e�<�YP��
~��(��z�O>�Ǐ?�����.��Y,k֜f��@��:�C����Ԑ5kN�z�I�=�+�7��>C�L��{a\��!r\��W��`h�Oݺ��iS�3:Ѱa%�Z�'-MƪU'����+g����?��<::�/��&/�`dd@�v5��������ܸ���>>W�={7NN6=:{�Қ6I h)J����ٺ5�C�nch�ϧ����k�NlaɎ�3}x�0���'�g�uժ6T�j�ر�x�&�ӧr�X�q��pp��ͭ&oߦ`h��T*��J%J%=z��W��z�`5��'E=�P(XY���C*�s��-Ǝm��k�]{�֭�X�bŊi��ի7����ן�㏽0 w�w�����\y�nak[�ٳ�d��m�|�?� -MƨQm5�M�'�oߦq�Zh����$'�ciiF�ڂF��[�Cu|E�@ ��� ���%::�)S<=���ۨ�D�����|���nn5Y�b nn5���0���Μ9�ٹ�J�c���Ed�v�¶m����P���}J�����@�f�i||��a�p���f{n�ft�^����!�+�~������""��{����dr���ҳ��L����I:�-S�ѹ@�K�{7/��t�\'Wמ<����*|<*�\��cǟ��.�֭��j��9}�!���Iɒf�^=�5tGɝ={6�?ִj�D	G*r��#���3vl;�us!%%�αv�iRR�<�9�ƹQ�T΂����s���^�ҥ>|�\��b��4lX�F�i���j���8/~~~l޼Y�f)H�n�4m�J�(DD�b��U
�*������ʘ3>,�����%S��J�T�4�����T�R�~�� M�D0r�Fbc��W �	�+��řp�^)����)���M2��R�֩M���S8p-�gwe̘�y.'2�����Wg==	u�ڱz�*T()��P�E==���c����V̑��q�9?�d͚���� ��,^|��+O�����ŽuN�]�h �{�ְ%�����*t�>�m�FӺu5bb���/�X��,
���C[�����b�P(y���.�dnU	���@�Z�*мyU&MjO�ƕ����}�v|||t�i+>>>j�dHU�v�?��S03�Q�D�ϱ�H�z�ה,����>>> :/z���E��f..���1[[KM�$�qD�V���H��)+�$��uk�8��g���< �#����
%w�Ѷ�,]�;w��';
���葞.���$�\ooIO�q��mf��Y\��ط,Yr��c�iev���xƎ����/����۷��MR[�l���?״*e�֭��ߟ;�Ō;�񹂩�_|ъ��[R��Ӿ��
��#0�	.<���'��'caaB����ט&M*��b_���?��Ζ-[4mF�����6Am�v�Y����Jbb*ӧ�����L�؞�S;�iA�!�7ANі~8!!���R��K���wyG��%��R��LΘ1�05-M�~�ٺ��|۠�T{�)�#6�m��s�4 �>IIit떳�-K���̈���rUOAp���`m]��'�|`"]E_ߜ!C�����}i���w��+�R9�n=�ҥ'����o�(UʜF��2Ń�M�P���H](��[�^0f�&���ضm4-[:i�$�@ �Z�r#Gn$-M������H*�s�x ��zH$sj��J2��?׼�II�'5U��5�N��щ ���:��}7h֬J�\��ߏ`˖K��K?LM�g�\�T�l�1~��(�{7�>�*��C�HC�P�f�:v������4�.�p��c.]z�t�L��4iR�Y��Ҵi�"�C t�R�ڵg��4n������VD�@ �)����ʕ���N��:�}���>��;`k[�ҥ�Q��	ŋ�`ff���ŋ�P��ߟ-,L177��̈/���o$�/:%z�ƾ��b���RS����o����o�݃��={�ϵ��"!!�	��C��    IDAT���,\�)�7״I�|�T�X�j0W�>姟�p��cn�xNz��r�,iڴ
����qc�\�X������[�p�1Ӧud�x7��-ٱu�%֯?˪U��]�����󛤲��N�QQ	��K����֖S����Nǎ�?z�#w�p!?�IZ�����+�[OJJ:�w��~}M�$Pffu�^}2�+7v�_�&4mZ;�R�6O j�ر�L�����M���H�z��6I ����'̚��)S<���E����=��122�����,��С�4j��Q���t�����O���Z1?�����o2m�vj׮��U��۫"�H>��*+��_���iڴr�c��%��TP0��SX��))�̟�o����ۈz�\�5�@�Ȯ��_����kF��@���L��A��h����w�?���kmW���DE�AOO��� J�r��K��u>z�ڵ���Nd���1S%��
��~?c�l���c�!x�2Y,=z�
�#�ܸ����իOu��.��L�����DA�{7�����k�aٲ~B���۷_0�>._~R��|u��E���$$�2d�66,_�_-�<=]Ʒ��e���$%}8��&���V*����k�	���x�:	�R���5�����F�.ًQQ����?cǶ��Khl�[ƌ�ĵk�X���V�4����X��$+W��l����O�zԨQNӦ	�Q(��^}�ŋѰ�۶��\9KM�%�A��ɪU�X��e�XЫWz��O͚b�^d2#F�'>>�&�-�CHH4^^g 022�C�Z��Հ6m��;;�:x'\d%�E/$�=��IK�������[���ak��cɒ�XX�2vl����/n�z��00�c���8;�ר=���]��=��+��w ���}��*�;��^�>��$�#��y���V�d�r*W.�)��ۗVI]9��Y�X�Y]���>t]V�d��?�����$����*'�ϻ�9�����>�]�}V�r�vu��EF�a�ĭ\����;��V*PzzLLHM���ڵ�Y���*Yӻw<=]qp�RY}yG��/}̆܌q*''}TN�����e\�m_����6��7{�v�~~�>�>�*��e>|�nbnnB�n.|�i}�4���>���N�on� y���:srL[Щ�-��o��X[�,{�\����;t�R7��#ٱ#��3;cl�9�h��@<=��ɆÇ�
�#�d5yϋ+��׾݇~/(X�R9 O�D�t��6]H�N?�~������!'�?7m�c�嵾_����]��yf�%������YMTs+��������k��U�E�vK���o���"(pލ�O�F�l�1�5[H�?��u��Ȅ|���qD���Eu�c9�U9��/V�\A��� ���"+W,p�%�L�R	oߦ�k�z����u����q���|�����U[W�ت�B���|��u��^����I�����V�Vc�Hd2s��e���L�������(�j��r���/*(� �eL�n�#(ȗo��KӦU�ի2��<�[�/cy���ש�n]~)-����������u�UW�֛7�|��^v�J��M��;O����-�w�ݻ/�?�y�|iܸ2�{7@&�``���17���}Ż�E���]P�?U���+��={��h�A~��S<<jiԖw�Ol�[֯?��է��+E�>IN���L���-eU����:%z��'P�L�<=���s�l]�._~�ѣwٶm�F��7o�9қk�BY�vH��
t3�:�+7E�f*�w^S*��d������?XѦMtX�q�:��c0�P��|�upT�v--;�~s˖�l�rQ�f�FF���f,d,\����ִjU �6�^+��Ϟ�*��x֬]̚��@��	��/^��OG��Ԫ�F�u��^�D���*�u�y�Έ		)���dI󏞯P(9t�6�5��9J�����eK'Z���2[s���Q�EZ��}�D���FZ�3V��i3
{�^# ��G��ӓdv�u�ؑ�|�D;:hmR�s�r��[�E�m')�&�6-Ri�� %Eʮ]W9w��;��g�03�Y˾}78q��G�{7N*�ʿ�� ��/Nc�C�ceA�_�F"��OTK��щ���!�3�m�-J���1���khh�T*�޾4Ri�J���u���#�}^�3�GL�[ ��sw�ڵP"#���r��mn�x���SUfgN9u��Go�jU֯���4�@.C�n.�6��p����	���!�+qq��W��t��B�R���߿�-�y4�1�dG����oT�J_i]�y�\0����T)^^C�Ǧ@cܹ�'�>&�H�'ԭkG�^���+�b*'s�|gw�&����nM�����*M-}ql�[�u�''||ƪ-SKVܿ|X�xL�]f�=\qv.����c^��n��{^�:#z��f����9:����T�R'��Y��,ZtOOWj׮�2;s�����n={�gɒ>��m�:�s���:�C{x7 U�Z�>}��'�(_��Z�̫�_A_��2�ca!� d�EU�cE�-����p�6l8G�N�����XY�,�@PP�'32�5�G��T���q2?㈺�Eu�=����Wu��MIIg�`/ ��G���!���XXӣG}z�p�a�J*	���3��{�ݽT� '�Lai[:�6���#��#G�f��e˖��|Ƕm�Ub_N�J�̞��m�.1{vW����E>��-��>���.�P(�J����KһwCz�p�jU�֥�����������(�?9�rz�rso4Ѯ>VVN��v�]e�ĭ�~��o�}Χ�6дI
���TY�8Y���_)�]�V-�E����qD�}@n�~�)KUcg^�ɭ-�yN+��:t=Ϟ���7�ҥ5' �{�711�s�:��Q��-�04T�0U����]��葐����>%K~�!�$44����������?eȐ��ٕR��Y��u#Fl��ݗl�0����^�@W�\��!CZ���J�z��H 5��d,]z�U�NҦM5v�Gٲ%4m�@ �� 0hPs<=]qu����G�T2e�6n�|����M@�Nޅh�đ�����QC��UX��&tJ���ףdI���{��]���Q�^�,�o�p���tƏwW��Y��AC��C"���'Q��m��+���5�_�&�6�d7��@�6W�\�_� ::�����V�G��I߾��۷����3�򢪾N��Lm�GS,Zt?��l�2J�I�����@�*,[F
:$z���/ɑ�q��<<je�711�?�8���
d����A���Z�*��5�R�>�yF >Ā%�7�n��		�,\�ǟ^�ݽ&>>c���ԴYA�D�.���[h�=����<�q����ӢEUM�S����ZtH�HA��R��*���y�9'f����u�\���m�`�?Y��,s��ҷo#-��`��\��~��'S��9zzz���͍��w133�����u��u�S04�᧟�бcm��X ��#G�0k�n
+V�O�i�$�@ �	v���ٻ�3�+={�״9�B�N�
�K��==���066�U�j�9��M2�W�d�趔(�q���"�+�;ח�1g�X�����է >��F�P��S�B��D�v�Ĥ��D���o�֭����Q��Jѱcm:v�M�F�����x�@ P��	̙��Ç�ЧOC������@ �#G�0y�6&Mj�5�I��O���̈%L133���ssc,,L033��Xg^�u��3		)H��N:��K��ղ<�r�I�1����$))��c7s��#V�L׮� ST��0�U+'Ν&=]��k�(^ܔ�O7cc�P�j���`�^��[�^p�����ڵ�)U��Zt�X�V��n��@ P=J��m��??%K��mۨ,Q�@�7ΜyȨQ�҂3:iڜL��]���==	��F��g"��z�����%���|�=��Q(����HNN���G,Z��?�bb���u��S;P���Zl��|�������g��gH�(���ʹs�9:W__g��l�0[��l�f�H$�����bϬY]x�$�Ços��v��!m�֠c�Z���T���@ e�<�fƌ�\���#Z1}z'LM�4m�@P���ű|�?e�X`k[+��-[�2e�ceU\x�
�̕+O:t=={�g�|OM���k���gIO���BIRRIIi@b����us+~aBgD���d ��g�<$=]��[���� �3f��j����X���L�޾�Z�)�t�X���w�$P*a��̝�=3և�������������7΍q�܈�|�ѣA9r��S��T*iڴ�_�`j�@z����OO�\uz��i3T¹s���%ajjD\�gΜa�B�][���H�b>�o��TΪU'Y���+���o2u�ک�.�@[y��u+�M���J�$s�1d����(V̐R����0��҈��)V̐r�̱�1���(�+�ח�����'����;/8p��5Y���֍�nnάZu*����Ipq����U��v���E}�b
j^�3�Ǜ7�Gv�G�ܡA�J�������y����ZVmN�|��Q�[�/��b5�=޼I�ȑ�<xSS#����1x���@}~��s�ww������������ٹB"1�d�.�}{����9���(��hcS�A��1hP3R9q���aѢ|���ֵ�@�����k�,�*UB*�ҧOM�Rd�T���M�7o�$ӧϊ�~c��Ew��#(G�GGoF&�U�qE������ܹG|��^�?�e������-(Z�{���3��fr9�{�J���$II2"#S �_���>"◂2]�/���S�xc�Ҟ������P�d�ד�q���W|��j6����Jo�F�*Q��1oߦe{�����ɓ;0yr{����={�<3;
b^(Q�H>'�Y�}�JP�J��o�W�B��˷�ن����ql��}��{���Vy|�M�.��׻�����}�l���y't������GH$Z����uq�o���a`���]I����J�2�:�H�r&L��ѣwX�r;�Vk}ii2Ν�ȑ;=z����8:ZөS:v�M�z�Y�k���c)AAa�t���C�P�㏽4��z�䋰�8��ߏ��M<<j��w�T�(<4�w4k���И��w�aQ��ǿC �қR�*J���XP��ۦXRv�4��$��ML11���Ę�1�����XP�(һ �af~�L����� S�=w��{�y�{�������v|��Ny,�-���س'���T�=�L&��ǎ�wBB<��j�
���"�O�ww+֯���*�JRS�ػ7��>A~~�͊�>V__SSC֮}�����G�hM���f
�����f���e��Oؿ�%��,շWT�1t�2^zi"�^S�Bɻ�n�/bx�0�~\�-�3��j **�;Չ�� W�ý	��ظ;���xy��\���D"!<܇�>�A�^m�k�=��
�,���?Ә93�]֫P(9q"���d��R��)��ܘq�<�0A����"'wi���yg��Y7���C�~F|��<=��U�P�U��ѿ�˖=�رn�K:�W^�¦M�n�� T��u�孷"�=;��Y����9t�4���b��S���`ii�رn���3r�6O@��2c��H�6�[�X�Ix\������))��ܼ7..����k.Ъ��K��f`l�]C�7�I���F��_�{w}��V\�1+WF�q�Q����}w�7�r����Fkll�� ::��+gr��~���Φ�����d�oO䯿Π�Ӓ��!4�#�k?�M[Ñ#���HP*��#x�ё��m|�a+WFkl�ⴴ�K	�d��06�Θ1I3ƭ͚�
�6*-���o)�ڍ��H�����u+��!&&��_����*�}6�'���4��U(�J22J8v,���,bbҩ�j�a��D�:�v��g�>c�R�$9��}�N�o�)������e�pgBB<;�[۾��ΔU���ۖu���l����/��T�D&���eKh�!!�xzZS]}O�ׯHz��颧���� 3f��+nF+���U��/��Ԑ��e�}��ɟ ��\1sKee=C�,���ǵ�	huu�>����b���1��r;���[	�����t�Ht��z�ƣ���O���~�|���fݺC���o,\8�%K�h�GAA%{�� G�f����ȑ΄�I?^zM�A�VU����,_����7H|H�H��'������!�(��,o���w'3q�K�F`m�G�a	�F�dr��
���R':��044`����[�f���>W__��=��|��]��_gWVVˁ�ؿ?���t��qs�d�XwBB���w��}Zrr3f|�����������r��'r�����0z�+!!��F��F�<oҤOHH�E�T�(��j��_>���5�O+���e�����q��k��_^^����[���y�o��]|��a�[�*C'����={-��ٰ�q\\�F�����ٽ;���9|X��V%:BBn��\]]#k��GF`j��'ݿ��s�m�����o�WYYOt�j&�?�8Mc��¤L� ����F���������d�mK &&]]\\,HN.D��r����.��:|��,��}n�DA������Z�k�>������A#�����ر,�;K\\.M��gȐ!�����V���Maa�z::��\�N��w��㸮D&�s�H��
$'�����Fh��G�`br��4��f���_��oϺu��kE]UU11��ݛ����j%�~�j�������z�~�/��SO���'��❀V$=RS	�OOk��_���͛���K�IM}G�ܨ�n`Ȑe<�t�5�M�FZZ1�g��O��l��8��y�YEE�w�*:�D__��cݙ<ٛ��N���<�΂�0b� ���/�kq�B11DE%�wo*UU��Y^� ���KL�(tMM��ߟ�֭�DG� �+
re��¤466��}e/"==],,z����L�3Q*�DE��l�6Ν���BY�0H�
]JUU�UII�dr��L�	�!Co�ttѢM���q�����`bғ?�q�FA�df��wo*��ر, p���Mg��N�'�#$ĝ��wn�|�fd���*as�x6	�Ș1z�qcݼ�
f���+�3r�6�ZhmZ���""�3��ק����ǿ���?������?��W_�Al����௿2�7oR�5_����9�xyy�v%�cG"G�dҭ�cǺ]Jtxгg�h>ԙ�<��ܹ���Ւu���Ly{hnVp�h&QQ)�ٓBaa%��}.M�+%0�Q��ZG.Wp��i�n�g��$��	HD��'{_�>�={-�q�\��]�f�\��tf'Nd�t�V���:՗%K�E��K(.����,u�##� u�����E�-[����5+�7ޘ*8v155��Ic߾S<�NEEvv���θqT]��ǣ����ν�e�h�����f��d�^U�������&��.H+�����̙_�źu�^q�L&G*}�_���y� Օ쀀�y�����{Z�֭�<��F�¤�Z5K뚞�;W�����ؑ��#g��M��w&MRUt�Dǽ��(aΜ/��C��[�a���4�ڽ[�$#��>}z�j�:z�K��-wJ�Tr�x6[�Ƴ}{��u����ǔ)>����D��O��3 X�h<���Bw0gϖ�|�v�Nf�0'�|s*R�����6�T*��,S'8��"?�<���xy٨���xO[**�x���x�q�Ԋ�@��r		yDG���)N�*�W/F��R�dϞ^x!�E�Ʒ��KKk�������ww+u����N\���"���#�|͌CY��+�k�9|�5����_����;9~�����N�k������X�`o�9Uk��*+�e׮$v�L���,�Lt���WZZ��EQQ%�|3M�tK99��ڕDTT
qq9��BX���w1K��)���֭�V��bAD�~�ۛ��2���={-O=5F�uw0ee�|��~�����S	v�tX�Ъ���IJ�'66���lN�����zz�솟��z�����	+�    IDAT�X%����*��RX�f?EEUH$�R�0//ۻ�@�P(IJ�W�IN.�{w}�w"$D՟��JT�	ӊ��o����ς�y뭈+���v�sg"��*���6�]Ə��w���)J�.��W_���oNe�����4�����;ٱ#����K��ý3�M$:�ACCO>���fժ�L���n[YY-��)DE%��gP(T�3!�ٳeDF��ٳe�ٙ�KD�����Oh���|���Ys #�����O"*p�PU����'8���hjj��̈��0t�#��xy�j�Q��uU1�7de����3��M�}�Rٷ�EEU��1f�;cǺ�z�~�����Ĥ�����++�KI�w�+�iE�cÆ#����{n��]q߄	��gϻ��P�?\�xG��~W'b2��g��Ȯ]I�Z5�)S|[�5hBii�v%�}{"��Y��э�w��}3ƭ�4��J�ro��7���k�Mn����Sm�ELc׮dL����Ԇ�0O�¤�RЈ��*�n���N��R���1��>DD���}ScwU��
6m:�GEq�BO>9���3�S�ͭ�ر,N�P%:Μ)��Ɍ!C	��!:��X�����3<��w��gȺu�]3��SE�����T��ёp�}N�*��m9'�\]�q�H&
�;ƍ�`�Xw�ݭ4��NH+�����7#y��p<H}{ee=R����1Ə�D�T�oo[>�t���&.\ϱcY�[7�#�[�U����jv�Lb���Ϧg�n�*:|v��W_��ҥ[�5+�w��G��R#�����3�ޝDtt
ee�88�c�D/Ə����A\y�LEE۷'������݃����~�o�����R�d��dV��Mv�9�������i� hBs�����ϾT͑EYY-ݺ���m{)��p��8�-47+X�� ~��������ਨ����t��;ELL5511�D��u'8؍�w��]�T��]ъ��M(��k:�:tF�9��N�̙R֮}���QSs��s�Gff�7?���]������ص+���9q"�^�	q端%8�M�UY�8����m_����),��/��Y�4A__��`W��]y�i�������ɬYs����?^U2b���5�_M�E�������С�t�ϸq��_�
rӒj�}�N��Q��0y�7���W��N�����ǳ9y2�c���GCC&&=2đF3d�#�޶b)thiiE<��&22�y��),X0���\��H��Y�VTz���.>�t/k�>Lx����_����%l�� >�_��~��;Z~YY-�f}Aee�6=���y�������'O�Ы������� W���$�y���ѯ���@��V��(!**�ݻ�IN.��Ѐ�`W&L�b�7���tb��xQ�޽�DFƱ cƸ�Kh��㫥:͊����#4ԃ�_����(u:���*bc�8~\����(A.W��Џ!C\�∓���4���L&��O���g����c�ʇ8��Ϲ��-{����=zVo�V$=�,����>�w�- $�]}��!o3c�/#%��q�>���uG�j��U��C_���Ï?>��M�m�XTT�Ν�'O�`dd@h�'�����+�Taa%s�|Iu���~֚��U�gO2�w�p�h&��#��0���P�͍5����dr~�=��[㉊J��E#F8�Ǆ	R��{h:D����f����8r�,������NU})t2������r������l
+��������*����H��
����c��M��U��7�Gyݡ�.4��_���ȴ����W�9p �s�D#S��iE���~d��X~��i�u ;�Ç/g��g���n$-����n{����̜�ff�l��8��u�1d����ؑȎ����bdԝ��=�<ٛѣ]D�CK��\d��o8y2��>z��S;o�[��j`��T��I���te���3a��	��4���B�ѣg���cǎD��/0x�~L��M���A�%$�b�nbb�>܉�^�H@� M�%ju�<����9�8�Mbb>/�01������;0 ;1u�Щ��\����n�!�������]9�{QQե&����W&/�Z}�ږ*����V��������f1LR�hE���7��/'ع�y|}UW{֯�����AJʻTT�1d��|���M��e�<��ܹ_��f����;T�}A�*ѱsgqqyu',̓I�D�C�57+X�l_}�O=5�W^���n�lpz�.^����DE%�Jee=..��Ʉ	^xy��U�oee=ݻ�+�D||��qlߞ@II5���S��v��;�u�:U����b��T�K/�1b� M�%tqr����bc����!..���s��Hpr2��Ϟ!C��� ��ZC&���ׇX�z ��:��3�"�H��$$������8u���=�1r� BC=;�s��mWii5����wo*�����	kƎu#4�__��N���.F.W�l��<��H���Z��x䑯��Na���psSM���_�T����X�b7?�x���7n���d��c�>ܙ�k�3��矿��H$>>c�W$:Ds����O��?1l�k�̥w�ѽ].Wp�XQQ�DE%SPP���	��K�0���@�ۚ�F�Tbm����Exyٶu��]��(!22��[���)�ѱ�:���*	��̙R>�0�;��a��+��
B{����ɓ9�*9���ϥ��CC|}�	P%8���i�/�`��d�-�FII5�橧� bb�ٷ/��ө���ֶ/!!���s�}N��G����#G2ٻWUe��SSCƌqc�Xw��\o���j���5 tt$�5�U��t�j��hE�c֬/��� 6�ll��ܬ���5^~y3ge��̟?��w�emߞ����S�����35:Uh~�y�oO`ǎD�Չ��pF�$]Xbb>�正[7=��f..���%'\J����VD��=	u',LJp���8�8q% AOO��K���#�7x���*���g��8�Ҋ��2a�T_�N�ɩ.$;�+WF��'qq���'0~����&��RIff'O�\���%3��B��c�����s`Ȑ��Xh}եе�<�˲e�8~<��S}�3�>��
8p@�\T�������3v�{�;&��(a��S��w��ǳ�H 0p cƸ�~E��͛��hя(��c}}]��X�z.AA��z	B+Њ��C}��&1�m��7�ĉl�LYş�ʑ#�,Y�'N�I߾�n���?̫��£��`���`��U�cG"۷'�����IO�¤���0b��Htj��u,X�))��Z5�	��Icrs+ؽ[Ur�D6ݺ�1z�aaRBC=�x���N>�� 2� �D���|��L��RJKkؾ=���8����۷���L��G@����+t>��\͖-�������ۀ����IL�WO{�DUUtﮏ��-�  @U�aj*��
]É٬Z�����pw���Ɍ��|rr�11�Ip�+���bb�9������Ig�^UeJUU�U���ۿ��N��Y�~����|4��2I�褴"��)'O搞������G{��c;��������t�}������/����iM���ؑ���$%�ӧO�K�o����d29o���~{��e��.�P^^Gtt
QQ�:t��fC�:&%,Lʌ���}�����ҿ�_��ޢ���UU5�kW��q9r�^��&e�T?F���
;����V�j�>~��VV&,Z4����ہ�frr��CUbc����Z[�! `��J{�Rq&t9�y�>����l����ŋM\� ��Ւ�cUMHv��Nr��'rط����"=��=��pAv�����0h�9_~��-��:�Hz��}DRR��#�H�:uNN愇{3{��<��]��J�T��;�Y�6�e���GG�K�99�ꊎ������>�Y�	wd�ƣ���/�����s:T�]M��k���4v�N���4jj.��-;�%K��`�(QJ������N%22���ttuu	q'"�c��}̯�y��u�^���;L߾�x�q̘1D�d
����"��)c��s��ϣ��}}]�R��<X5���E�4Y��N�P�n�!��"���*$���e�g�l(��}5f���x����n�==]tu%,_�f�l�Ȅ֠I�q�>�ԩ"

>���"��z�6m�`��ǯ�<�\��/n�_N��'���~�6�3'����ؾ=���B���ń	^��{3l�Ht����\���CC֯�'��W���������ͱW�-^MGG�ر�Z5��4�m+MM�8��֭�DG���,gԨAL��GX�CCM�(h@yy_|q�o���^�����!̝;L����Y���%�<��M%..��g�P(�������{|}�JmE�U���ػ7�u��Gs�}��\y�!�5�K�r���[Y��MM�[<R�D�$,̋�?�!�;	����pA�N9��B���ʄ��`Æ��}�L&�'�%&&�u��1v�[�Ė�Sζm�DGjj!���L� eɒ)���KÄ���ߞ���?=�&������:}}]RSn�� �����>_}������v������n�g׮$��.8�7ߜJx�7}�ܼ����Ν�e͚|��aX�8�G�!fH:���j����I���|�044��ۖ�0)������cff��pA���ϳo_*۶%p�D6r�	������c	���w'�F�@�R	{�����ڵ���y��z��􈍍e�С����P\��!���10HCC"={zS]��ϒ`b2���d����0������ŋ�\�x�ŋ�ɻ��f����f^}�~��O=5��_�(��P5���{��-n���A�T�A��sa455�q�ڡo�	���kǔ)��WD�x�VZZ��{�~8B��=x�1̝;L$;�;r�BII�����ɓ�W��#a� |}���W��pv6�:��_�w�}W�ah1	��ϢP��ܬ�oߞ<������/H��3l���=�R��%P*%��=�N�n~QMh?����s���5���� ����U�zಟ�]��F�v<Vs3��Dbɻ��ANNv��O�u���g0�W_��'����v�����Nx�j�&��Y�l��5
f͚Նv~7ndǎ?8s�;�i:AÊ��X�� 7�o_C^=�ٳ�C
�[R*��={���\r9y2���"����o���=?<??{||��P9-������>6l�t(Zi��9���:t��d�Xw���%�affL}}%���J]��]�=t��M=t��]]�uӥ{w]��5�_�M~B�ٳg��}����<����2�.��?��tB2c���mY�p=���z�F�v�tX���@�^��H044@"������G5&����D��Qwtt$U�e��M[��i�4g �Ɉ��	�.����ի��q�Q�̌y��f�*zv7TUՠ���j:�Guuݺ�!��8��������7S��M�&��m$22��<�6=��P:{{S��V��f�aÆ�X  DFF^�vq"Z��Ւݻ���[�={-�>ʢE�df��Q̟?ꮞ�a���!�����Z��͛c����;�<�C��Whjj&%����<����%+K5���C?���y��0|}����ۏ �"]�N?� ���-׫��W�!0p K��ʱcY|��l,-M4� Z '��U����/'��2�����ɪ@s��3gJHH�#11���|�Ҋ������׎�S}��U���۷k�AچHzB1g�}�������!~8�	��K�N*;��~��_=���)+VL��,'wQJ����r�IH�#!!���B.\h�G�nxzZ�����c��C�.;K� �оD�C�ww+���曑̛���so�9�K��.½��,��O���C?V���ԩ~"���U]V���^Ss}}]�ܬ��塇���c�����>A�IA�bz��Ɗ�	
r�~���,>�|.nnV��K�H$w4�Lk/��Jkk� h���<֬9��]I89��j�l�N�EGG\��v���_��HJʧ��	NN�x{�扏�=V�i��!������w��X엻�U�]�-��vv;�n���{����m�W
������\Ann�D/|}�x��L���W_�����D�q;�����>�-�)t]11�������L||��⋇�8�K$;�T]]#����窓�����3��ǎ����C*���
�=�|_,�˭gӦc,Z����Gᇟ���C��������_��{I*�j�w�Nb�4���.��҄͛�b���,[���{S�������th� hPs��;����ZHP�+�7?ňΚMhE����T���HH�'11���R
%���xy���CC������N4����,��o�⫯���ʄ�Ӈ�ˠA�Nho���V��R��r���{�叻��;��hy^�2�f�W�~��o�A�tt$<�L�G���;vo�}?3f�th�VK��z%���w���=��������2/���H�y��\��ĦM��]CQQ%�'���'3���th�=jll&=����|��HL�'=�X=����-��{��+���3|	����n���w�}���s�+�W�/_����&��FGGB��z\�����^��O>���ٜ���:կ�.�]=D���W��=��|YWo;�Z�ݼ�����U1�vܷ�*I��%<x�����~�	��w�N�1�j9�Йy{۲g�bV����śؽ;�>�N��F��S���[=�^lng�w��}JJ�Y��?�p���fzhaoo��Є�p�B���$'��\@RR>gΔ"��12ꎻ���7�'�3�����n���9k����پ�5�T��� df�����Y�|'>>�L�6��poLM�j�7JT]}������z����?�(�r/�H[ns7����빑6�r�D�����D��Z�N�)BWe`�ǒ%S?ޓg��Hp����?���:��}X��}m�е%&���1�ؑH߾�x�� ��&�1t"��/%8
�_��e��
��{��e���.���c��R%8D?A[����vm���u7모0`���6���)(���}J��	���|��
X����l��u�]���*��}���6	p�	��Z^{j��ǝ&���h��NM�.�m�G��}�����O|�Ν�,[����- �+ؽ;����w��F*�ᣏb�T_��u5�p55HJR��zq䓓S�B�����Ԇ�P/C*��:�p����v�J�֎��i#��V]fGu�C�
%�:Q������Ъ����uu��v��^�Nb����*���o�j��;��f�6�Jk�ST�]���+VLg�D/^~y�G��[oE0}z��C�.TTԱi�1���0�����ɯ�������M�����+�7���ͭ ����Ԇ�?<=��Jm����fngXi��Ek_5��r6l�Ъ�쨖/��W_�~��H$tu%(J�������g����]S@wS!Җ�ެ/H[��ڤ�ǝ<�-�l���N��C�
��\9p�%�{o��ȯ��dŊi�ى+�7#��
Ell���Ů]I��ٍ��x�ё�
�)-�Q��HNVUq�J���� ��0}��R�R�͍5� tLw�����;*q\�:$���A&S �Z3mZ �ᾘ�����mS���o���������m�������˓Wϔr�$��&n��;]���wA�
z�2`ٲ�����61f�
^~y"�=6]]M��!�h��{і;�[�D
�Km�E~��$�~�'%������Ә:՗���5^�VXXyixJ�:�QVV���)R�?<��OO�n�']���n����������u�.�_n]����dr�ϴiDD��Z��f�Э���Sit����Ͽ�m�-�����Zqߎ6�r��/��F?�l�wý�S49�������}��w��Ndd�?OO1���ܨ���~���nw�w�>�s:y2�MS��_    IDAT�b���`�T_>�l�x�j�L&'=��S��8u����"RR
��j@GG��C?��ly��`�R��l06���ӹY��vw�}��ｓ��f�,�׷�P(��՚����<��nnVm���iR7�a��>�u�i�X�{[o��[4A5�����ˢE�4ɛ�^�̄	����'�vAЀ��j~��?�Kffnn����$�� ���k:�.�����tUR#-����BΞ-C&�ӽ�>..xz�&���k4� �֚4ɛ��ZfϾ����t�z��u���͆�<xP=�v��bAd��l�r�w��ƶm	��z8ӧt�1���f_������ٳ'�͛c����Ȩ;������s���txZ��YAff��z#%����"���޸�[��sυ��f��c1P����v.��v���j�u��H_�Iz�n_AڏD"a�� ��<y��ݼ��Ol�p����ѥ���zg'v�]�B���ѳl�϶m	��^$(ȅ5k�2~�'ݺu�]z�PU�@jj�N������dr��uqv6��Ӛ� W<=�pw��o�^�[4n��DJJ���3���;;S��%$���͈�cGH� �3c����̜9�W_���?fΜ�x�	�$@�R��ĉ�mK`ǎJKk�����Cx�?��{k:�NO�P��S~ihJ���!*-������n���N,X0ww+�������p��1-X������텝�)NNf�ۛbk�J��ۛbnn,*DAhS"�����{2a��xz���yxX��n�pA���f�֧ټ�8ｷ�_����1o�Hq� �I�T��T�֭qlۖ@QQnnV<��H�L������C�jk/��^|EGZZ1.4���À����ᇇ_�?[�Ē ܡ3���/'hn�{�����9����|tuuin��P������ҳg7���2�BSa���Dң��<ؑ��B�m����"zz:89��d�RU"D*���H4�:�DC�<ٛի��b�.���/^~y"S����9�p2��Ç3ٳ'���T���pr2c�̡���0h���C�Td29����9SJZZ1%����[�R��ظ������1{v ��ָ�Zb` ��^y{���/'�{�\�D.o��6�LNu���M�.J��ۙ����K# �ռ��
��HN. 5��U��QQQ�D"�����F�qw����Xï@nO�^���D�̹�+v�}�W_��[oݏ�����������iDE%s�`:uu�xy�0w�0ƍ�h�i��Is����s��s�t)�O�����hnV���ˀ�qq�`�� ��U�7ll�h:tA�Z>>�WTy܌��J��Fs��tuE_AZ��K�.m�8�Ts�zzͷ~�M�/�УG�=�ìYw�H$88������>��KJ�Չ���B����+���Y��a�����V��X��B�em݇O?�ł�y�H�L��ɓ�y�	h���n��ٳ����tږ-[4B��T*IO/���tbb�9v,��Ýy��Ɍ�Jq=r�������O���Y�L&GWW;;S��,�4�WW�`�@3��v�������T@RR�-����Q�������4Ȃٳ7�q�Fd2Y;F�ulٲ�����v�y�h;�(��D*))���G.��[p���Q����TW0`@���pv�B"��B#��z��_����e���I#������xױΝ;����;~^UU��{�j���|cc3���hv�
���J����]�)meϞ�{o'��e������=
^}�U2335F��������5F�QQQ��g���ĤSVVK��F�9�q�<	vC/�T*��?OFFɥ����3�\�(CGG��m_����WWK�`� s1{� ����r��
�蒒�j@WW�����!66�����}����{��� "�W=�u���|�����R���=�J�v��]o;�&����3lػ���3!|��nv�|__;��j9r9����z���O�9r�,C�:�쳡��⫸s-e�iiE�����Ww������������@�q�B�d��x>�x������y��q�ٙj:4A�'M?���Ù�Ĥ��Z���C�:2z��G���a%z� EEU�>]�����P%7��Ull���l���j�WWK����ٳ��#��A�T��]�Nl�Tr��\@OOggs�R��l�����Z��|�_����dsi�2o�(^xa���xT���I���:��%�ٙ2u�/[�g��a<��8 ֬9�G��?^������;�ŧ��%&&__;�}6��P�u [Uՠ�L��V̩SE�9SʅMH$��d..��ߖ`ggs1�����r��z��+�),�dƌ!<�L�o/t�����fs��Y�$))�L���9#Fb�7�o`�>Q/+�%#C�L����3%��\�ܼ7..�}Y2h�����v�P(��:wYr#���Bjk/����������^s7�y�bY�x
���C䀀���4\]-��U	� �hE�C&�co����X[��а;�O��m�3 455��Ԛ/�x�U��ǧ��e��T\]-x�`""�:��a�BI^^�e%ê��gΔ��Ԍ����}qs���Qt:9�w��$h��f?�|�O>�Kqq>��O���yz~]CUU'N�p��Y�=KRR>��
� 0БaÜ:t`�k:�ܬ���<gΨ�+gϞSϞRU� ������������{��p�е��
23ˮ��HI)���}}]\]-��//�ܬ�xf�ӧK
z S�^��V<�ߡ.
��uhE����%�w����g�	ᩧ�'9y&&���={Rx�u���:Ա�֛�VĚ5ٶ-����X�0�Y�;M�^s����r�Ӌ�	������!�����Qw�8�ggs���pt4�4�Q�<d29[������}���|2�U߳�p��r�O�p�d.'Nd��ٳ� 4ȜaÜH`�@���=�����,��ٲ+�-� ++4���gg���ps����P��B�SW�Hzz))E����ZHFF	.4ѭ���V��T�Jp���.�BI@�ی5��K���XTn	��9Z����y�aÜػ�'O����k���s�2��YQf�����:����Ӻ�悂J��2���ҭ����0��M�~�� O&�s�l�:	r��� ��ٲ��''3,-M4���)J��K���r�X��v��_c	���{WZTT��G\\.'O��K]]#�������g����;���H�PRTTEVV��edf����Jn��TЭ�ޥ�|s���� t ������������[�R��ظ���xxX��f�TjàAb�?A��Iz����C���c$$���0�+W�T?&#����x�i̚�&qTU5��7��7����ȴi,X0gg�6Y_{k�6���9+�gΔ��YFe�jJ_CC�K��A��������r�d�~���d��L�?> �	�������|�WRR>�H$���o��������]]M�����j��*#;�gϞ#'����sdg���Q5�{߾�pv6��3�ֶ�V�M�3���9SJJJ!�Nr�T1))TU5�{�yxX��a���5����Q� ]��$=&N\����}w��~{��Gϲ~�_�Žy���%K~#22�Ç_k�&i/���X������.gԨA̟?��`W��R}�|��r�+���������!�0�ߥ��0�vv�"!"�TNN9k�����'P(�L��Ü9�����thBW]�@JJ��y$%������b���//[��U_�T�Q]�@VV9YYede����(';����F��z0`@?���hv�g3�UA茪�ԕ��"N�.A&�c`����%����$����h,�p�Iz̘�9vv�DFƱtiR���ľ}/��n�~\UUÇ/gƌ �xcj�ǥP(9x0����w:̀��7oӧt��c�����[�srT���j����ں�U	UR��ޔn����jj.��o'��#����nŜ9�x�Q���57+��*#=�X=�wZZ1����j����FK���A�ܹs��斓�[ANN99������Uxݺ���В��Nl8:��ܼ��_� J����
�gWJ�*����ejj���pw����
''s��Dŕ ­hM�c�����J�ͭ�����S��y�������^��o���7����_�ѱ�Ř�Q��_��/��D__�Y����#����n1t4������/����2v\GG���	��H�88���ޔ=��T�]]\\.?�p�m�����t��Z���zuYwZ�j���%466������f��Z��a���V���ef��<UR����{}}#�Jl�ۛboo���kIpX[��	A� *+�IK+VOᜑQBZZ�����a��~��[��is�zò�~~	� tZ��x�����V`nnLee=?���g��@QQ?���+�ܬ`�����߈M��h�X++�ٰ�(�|�'��Ռ��ܹ�3�M�^��&D���i�t��7�ֶ/66}�����N�Y:�������	~��())���1i��� ����d29����:UDZZ��E��� ��������..��9_EE���),�$/�%��JjV�H������臃CK�CUgi�[l�Ё��7r�L)iiE�%dd�?�LLz��j�����V�&��b� B�Қ�Ǌ�ٻ7�)S|�����ƾ�o����sIM}��n�Ǐg��>�)S|5ss�������0���¢7�f2{v����Bcc399���UPPp������W^�~^�T�����	�>b茖��:Gdd۶%p�t	VV&L��Cx�/��v�O�����ӋIM-$-MU�q�L)2�}}]\\,ԉ��$Gg�*���^����Y�R������&@5��¢7vv}��UrCU�&zlBǣJΪf�k�:KO/&/�<J���=���l����e_�XO��hM���/�������y��̙��p�	o�7��G	�^�E�6��￿��O99����~�)���BC=�;w�F�hm�ӶTW�x�IEnn������<55�~�33c��TI++,-{cm���XX�`f�9N��k���m[<[�Ɠ�S��Mƌq#8؍#��L_�����Ξ=�n�ܒ���荻���R\]-;��O��
��k)(8OQQ5EEUW|�VRW��ҒԸ<�zy����I�}����)J��*.�RLFF1YY���YG����X�榪�h�9E�	� h��$=�l9�K/mf���1b9{�,F*�aҤ�H�6��޴k�s�|=#G���ҥ��ZMM��ڕ����ȑ��ۛ2}��O�ں������WT���NNJJ�))��ܹZ�c��u��4�¢�:)bii���	�潱�1�_?#14��KL�'::���IJ�GWW�����>'��s�gOQR�Z*+��ͭPOk��թ��g��C5��L.M�j������xxXu�j��%�QEq�ꫠ����j���)(8Ϲs���
 ��t03SU��$SERC:���j��U-_gΔ��ЄD"�ή/�����2h�NN79+�ЕiM����4������� ���ʕ3y�>�`7�7���7�������3QQ����#8s�����'9���C�>}�'{�+�m�����bU������j���)*R�\TT͹s5(�������cm�K��W$H�̌���33#��{h��	�����:t�cǲ��)G__//[|}������G���G�47+(*�$7�B�T���*7���� �+�NN�89�]�2g�@�k�����JKk(+�����s�j))�������*
+)+���Y����ա#ll����66}����B�� �Τ���ӧK��QLUU�"����2�n� �$A�D�&鑐��ĉ+9z�uy�kƍ���W&�ǤI+�����R�dʔO�Htغ��y�#������l9Ξ=)���2~�'3fa�pgQ2�!2��s�j),��"A�r����&PͮЯ�!��DH�~F�~6T'FTߍ������#G�r�x		���"��16�Tjs�WU���l�%�7uu�URT��n(*RU8W��l�Tlw��N5c���߳��ٙbmݧ]�T���?_Oyy��U�D��	�Z��j(-����Y�����133��\�ea��R�+������R:!�B�V��YFff)�O_9��ظ���h�w77K�����A�{�5I���r�{�ݻ�f��r_}�(J���g�Û��?���&m��I�^�Qf��%e" ��8AE������U
zq���((��Q�2eʞe���I3���H)t7i���z�<��~�9�����9��ӧ�ży�*=���T��O��)}y�uSP��֭g�~�q�<��� ��1cbйs���Gw0���-ANNrr���U���bde�>U��-FFF!rs���[\! qq���
x{�B�� y�}7xx����
<<dv�K�Ht�2\����gSp��-\����W�-�`=慰0o��y�/e0�P4�O�u�2��!#Ci��LO/,��f7������r����|��f��pxy��@��#/��<�0��c~��[���"�c����\]]����;��u���~~Pp��j��P�ڵ���n�C΀ E��3_�k�6mL3�XT���Q9L�QTT����X��i�8��_~9�� ^}uΜ���;�Y��o��	?�|�o6�~BB6n<��O"99>5�+F����P{�����$;��itnn�% 1_����� �%6� ���������C�����\y�W����r%7nd���\ܼ���S�\s�J��	����Z
xy����>>n��v+�f������%((P!?���*�竐�[���B����5;����]R>��4���t#0����
�hp��ӕ��@�R��B�M�TW�\A��=���f.."xy�������94M!��SЉPA���lsa䔔<F�DB��y#** ��~h��mۚ�յ��zDDT�Ä ��,�1f�^�k�ރD"ƞ=���?����o"(ȣ�s��J1`�{<����I�<�;w.[���o��ERR�ý1jT7��]�2 qDEE�((PY.vM_U��*��章��+�#
,!�B!���nn.��\ �9C.������X��B&s�T*����r)�Rg�d�-z���p��qSS�Sl���Vk+���.���;
)�rI�� ��"�������zF��j�V�RiP\��RYj��q;�L��L3�L_MA���^^���C$r�l٬��+�O�T���Ci���:(�jh4�㊊J���QR�AI��EE�P�u�hLǖ��T��z߀)�0�o)
�徇��ϙ//7����3"j�F#RS��`�
�\�ʕ�� d2g�ic
4�5�ڵ@D����C�ݻ��>;��G���bǎ
�V�N����?�G����l9�g�����<bc#o�Vv�B*�n=��[� ))��^92�wD�ޑ�C��S��B������B5��K�Ri�Ri�T�QR��Z�-?O�Jc��Pww�ŻTj
L��L�L��P`	F��E�JM�»�:[~.
��b���Sz��..��s77	��
���,�ck�3�єUzQnVXh*f���R�f��Z�T颢RF��P\\
��%%Z��Zh���~�����T��Q�ӣ�DW�w忆�B!��+e�FXv�$S��������.pv�������Eww)�Rqy�!+�dP($�Dl��BDM�NW�7�q�����իHH0=V�L��}|�,���rpW;""��
=�Y��û���G۶���w�cҤ^ ���^�R�u�fU�ƤIː�W���_t��u/���_�b׮��O�����k�A�:`Р�������ʠRiPX��$%%��O�uP��(*R�_� ����̲d��TwGx`��`�������?z�"�D�Ż������J���,�\.�X�77I�q"��R�D����El�c�a��n��g�TF�ѣ�T��"�%1jp�I��U��c �
K�$1$��9�""�/�ш��Bܸ����l�K|��    IDAT�a�%$d���\��89	�e��Ѻ��eY
QC8T�1i�2��y���'bĈѳg+,\8 ���'��?�����]ϙ���!C��믏O�5��Ezz~��������PR�A�6~<��1�1Ou'jjT*-t:Ӆ{a��2󡸸�}�ۗj��~�_�\Za7'�B
� prr��V�DDMQnn1����]!�HḺ̨�˥���E�V>���KS�7قC����'GV� СC���,�� �o_<F��^e�[��gc���1"ڡ�Nz`����>�/t�2;v��]�޽�����pq�[�0���
�zE�G�xx��jLK]L�]���}��ƍl$%� !�Tg�t?�RcH*uFD�Z��Ő!�k�y{���QK�P3=�z�>|۷��+�����oY^�8�sxy�a���ն���q�}�#4�k�<m�a7	�����k8~<�uׯg ��УGz��D���m��-�� 11II�HJ�ER��~bb�e(��	aa��V�|��@E��rDDD��P3=����* �o���bde��� 0bDW���Vh4�j��;;���M�رK�a�qL�гQ�oO���8�'&N4�ׂ����O±c7�~�qh�z����K��
��0!DDD�IFF�%�HN6��9�A��"��y!"�117���MAGH��C�>#""��P3=�l9��_����QX�Fǎ�c͚�1hP{ @f����b�Lޥ��^}#6m:���ǧeO��j�8s�&ΜI���p��-$$d��� �B�.]B�Ν�����������Z=n��Grr.n�4�̡Fbb�������¼Ѫ�""|Ъ��ýዠ �[NDD͞C��_����ܹ���㆘�x�x���cƎ]��`O|���+)�`РE��	���3l9�fI���ҥ��$�Υ�ڵL�tepw��cǠ�n�h�>��E)՟�hDV��<��Crr.RR����Y���'����e�F�V���0�Z�Zf�9*[�" de)���q�rz�cF��ŋ�C���X%����O�ԩ_`��X�g���9�ɜѣG+�����V�G||:ΝK���8>��GI�B� >��)��t����)KDDd-Jei� �t?��~�e������^�F��6�3�ý��P�jw�#""rtz���z�/���\ᘑ#��?�ٌ}�.cذ�C���c�x�p�=�!�Km2vG��,B׮���5���hDrr..^LE||:��Ӱn�1����h4B.��S� �m�v�ж�?����9��Bn��ǭ[�HI�í[yHI�CjjRR�o**
�ﯰݺ�[{��O�¡DDDUp��C.�@"#3Ӵmmtt(��rJKu�H� �� bb"�m۹Z� �p��Ž����|��$���Q	�>9������R�ǧ��%Sr�J�n=k�#O���!�h��QQh��!!��㎈�����"���W2n�2��-C�lՐ/{��v	�DX�7�ý�Y��T"""�����@v�i�����\�����p�1�FuŒ%;�ӕA,v��M�~{f�Z�1cbЯ_[���%qw��W�H��Y����b\����׳p�j�]���ݗ,a�L�l	Aڵ��	���+����teHO/@zz!n��CZZA���<�̍�R ��I�� ��=�N�� $ĳ���P���Ȇ�_X??9��L����P(d8{6�B�1rd4.܂�bȐ�j���aӦSx���㏗!�� ��x{��o�6�۷M��U�v-W�f���L\����Gp�V>�F#��Eh��m��WC"#}kn�^o@V�ii�HK+DzzRS�V����� +��Z���"y $�������@X�i�Fh��w����N0�pGFF! Ӳ�.]Bp�\J�c��=ѽ{~��L�C x�݇1p�b���v��?Yu�T3�BvW�T������0���̐�~:���<�� 	�eْ/<�ޖ���Q����0���.�`����7����.BY�  	��'Gp�'��<ЧOky 8����`*""�&�C9.\H�<���޽��:�����waѢ	��R����o>�W^ـѣ��{�0����O&sFtt(��C+<���q�z�_�BRR��sq�jv���B�'t�
����{�� 1�""�桸X���ddZn��J���ff���#'�z�)�
���#$�^t���
��	񂯯;�N5c����A|��n|��9� `��3x���p��{�b� ��Y��؅�꫙x��.�n�h4bҤ���-��t�fJ�ї!9HL4}MJ�ERRRS�ӕ0�s�{v�O�p���5��YY��"3S���B���h(��V �Jk9G"# @9=��/GP��k@�AA������q"""�p3=��=��V ���д�E�7���4���]���_��}�`Ӧ�u
=/����{K���_��o�l��E��� DE���^o��[yHN6� �ێ瑘��F �J�ፐ�ۦ:+��?���jA�T#3S���bdd"'���qrr���nz�\�0��qG`�~~r�k�{�mk	4= �L="""ࠡ��!��B�s�nV= `����_?�����Z��W_���ފ�C;�K�k��#�Hh��u���HL��͛�HN�Ejj>�^����W��V �������oE<�ݙy��ۭ���M��ꐕ�DvvQ�0#+�h��!=���Ŗ �b'x{���_??9����5>>n
򄯯;��<������M����vnyKZZz�X��[�"66 0i�2y���T8V�T#:�M|��$�ߣN��FL��9rsK�cǋ�j� �~.���*ƻu+�r?55YYb)��-��̕�CB��@`��9WW;�#"j��zrs���W���b��Y��� /���J�V8���>>��������nP���p������//W;�C"""rdw���/�H$Djj�%�Ş=��:V.�bР�ش�d�C�@�%K�`Ȑ�X�h�����>5s� ��r��˫,t����C�����֭��A<}�&RS�QR��/�:�_���������� ��B��_oo7.�!�����B���dg+-�F^^	���~��[����
��N��r���+|}�����hOK������KDDD�d8\���$D@��n�[������{�Vk�ڞt��<�����)��Oݖ��za��1x�>�z�lU�I��9;�,�g�RX�BZZ!23��mZ�n^�~�rrrL��*��
�/B|}M�p���9����K�����/(0���S�����y�s%w��0����r+���.]B,�O������w�!�K��n�������B 	�Bjj��qtt(���x1=zT&���D��[Oc���u�kʔ>ؾ�<��]�?�x2�s�'�@��A���C��j��h��Ha�k瓒��];���
//Y�WWxz�o2xx�n{�tY_q�EEj�QTTj�zg�a����w�q�
U�DY���=ЩS���i�WooS����DDD��2��ĭ[y�������v�ɓ�w�R�3�O�+� ��ߟ�A�᭷~���o�؉���ET^ĳ�c��%!/����yy%HN�ũSɖ�n��0f��b�tAe��2�&�?vw���݅T��#�JS`a�ZTT
�R]~���ߡ���w�֒H�P(���Yn��r�kP!��=���t��5;9l�����
���F��ɤJ�;6Ӧ}���\��{׹?9�{of�^��ûT������R��R�m�_��Z}y b�>o�B��Wby��W����
�WV��]WW�� �t��C77	��Lϛ�+�
Ǚ�sJ=Y�F��J��RY��T*�j

TP���7
Ֆ�%%�Z^+**Eq�*�j���~�r	�ݥ���I,��x����U��Z^7?���DDDD��U{VX� �z���_�Y��������6m:�^V�>G��m����aϞ����=gg����W���ш���l�'�����EE˧�EE���V"1�|Y��5JJJ��*m����:C&s�T*������DN��%�E�ɜ!����"���"���I��2�3�b'��R89	-�w���ơ�PRRZ>k�z}JJ4�h�(-�A��B�գ��ee��ee�*��@�-�p�^_f�9,+��g0-+�JŐɜ��&�\.�Tj�y		񄻻��g�r���.�ɜ��.��u� C 4�w������ⰡGa�
���������	��ooEZZ��<*/	��ñX��8��Z�?V-�!C��K/����~�����/�VkQ\�)JL�LuL�Z�EQ�)Q*���ʠRi��Q�F_�Z��J�ՖY>����j����~5*R���I��$ ��:C$2�H!�:���t���Ȳ��� ��1��E��S]f��C��0���T�+�� ��:���]F�6� �Ri-�������R˲s�F#PXh*�i0��ڴ:b�d2H$��������B!<<d
���X�D\>�Hb	�n.X������19l� �����
  t�
�H�����C��:g^X�|���>}Z׫_�B��?~�'/úuG1eJ���	�L*5}����n����R���A�,�V��Z��\���+�/�M��k,��sL���:h4zh4z(���%�Y��eeW}�_Zj��P[������pu�T��\.�PXy���"��>�D"��<2��e���ii`��#�"spt{�#
��.)��%2�;��=<�
��c������ńR�3:v�ɓI��:"::?��W�C ���6�={�|s3M�ےQ��M�\�FDDDD�����-����$���Wx�W�VU3�I�z��_Ϣ�DӠ�_~��n������DDDDDDDd[z �mk+����p!���sƎ��NW�_=۠��b'|��4�ǧ㣏v5�-"""""""��=�¼p�fn��bb¡ӕ����J���a�����ǿ��6~x���������_7�ՍÆ�Z�"11��s��^��sǩS�� 0qb/;vII9US[ӧ����0g�(��O """""""�q��#"§��W��j�z��E��_��7x� ~8Zm^z���GDDDDDDD�簡G�V�P*���-��|llD�����?�?�t������r�g�M����jա�GDDDDDDD�����i��;g{�Ɔ#+��ɹ�� �8�'RR�p��5���o�6�7o,،K�Ҭ�&U�aC��@\\Dw�����D"���h۶��ٳ֬9j��̝;���5kT*���%""""""��9l�!Ъ��]3=��E��#�_������b۶s��)����rr�Ϧ!/�����U�$""""""��9l� aa޸q#���﹧M���ȑ]��&�?��x���裩X��86n<i�v��������nz�i���wp���HI�CJJ^��J$bL����*M�#f��W_݀��,��KDDDDDDD9t�捄��gz�ĄC"�8�cڴ{�������Xu\��6��੧��Z��DDDDDDD��СGd��J5

T�7��8z4���[��ý���w����b'|�ţ��*«�n�j�DDDDDDDd�СGD�/ T:ۣoߚ�z �?���q�V[P�>�t6m:�ի�����AApvUQףM�u= `��.��t����fqqQx�����o�ٳ)Vo��������%s��C( "���w����=�Vu=�b'L��k��^o��_xa(��o�'����%Vo���������r�� �ý��x�Ls]�#Gj^�2m�=��,��ݗ�>>�@�O?��@���ު;��dzDF�V��0��8r��b� ꅁ�[������_}�(��?�e�>�������Z�=Z��õk���ַo��z ���}�o�e$%U�4Ttt(�~{>�hvIDDDDDDD-�Ç���C�,�t�����kU� �¼�b�[�iͤI��쳫q���uH���������>�h�> p�J�]���N��#�V��P(�O��?��Rm�q����x�k�G]���f�9:�=�r)�� п;����Z�5iR/89	m�}��X�+f��D�9sXؔ��������>� �v��=l���B�ǧ�؎��y�V���&�ך�����g��?��vج"""""""G�"B��� \�Zy�ѩS0||ܰ��Z���c���Y��;�[s�w��-�M�����[�ش/"""""""G�"B����!
���]�U[���2�#���5�X�	z��'���!>>���9�z�k��bRS�+}}Р�8z4j��V�=�d��R�9�J��ߣѣGf�\���b��GDDDDDD�(ZL�T�� ���ռ� ����;㫯�[m�Uqrb���
�1ct�2��IDDDDDD�ZD���.Ap�'._������:u
�u]�4�c��S��TZk�U��t�ڵO#11�歃��]�������j�"B h��׮eV������� c������V���j�/����[�`Ѣm��'Qs�bB����\� �w@BBRR�j՞X�3���ՇPZ���0�կ_[|��,]�7�l�>���������z�k��W3�\�\�={�k�����B��cݺc�f�ƍ�ų�Ƽy�j]���������%jQ��J��r&�X섾}�֩����+y��-���`���h���x��n�5k��r�_""""""�����.q8�=�V�Rf���L%6mj��&� |0	��ޘ:�neKDDDDDDT�z��� 4ԫƺEE�8y2���(0~|O|������D"ƪUO  f�X�Z�h}5-&� L�=�^�:�	�D�6~ػ���� �s����ع�BC�X'��nX��i$'�b���PV�xKl���������zt�����j�����ֵ Ъ�/F�ꆥK�h���%"��V=���b�ܵUj%""""""jiZT�ѹs0�^̀V���a�:�T��ԩ�9s�������Ն��bb���O`��3x����""""""���E�]��@�+åKiUӧOk��K�s��:�ݩS0j��Kw7t��ү_[|��|��|��~����������)iQ�Gx�7
Ο�U�1b���;�^�cΜ�p��U�>}�!ì�q�b�`�CX�`6nl��d���������zt��s�= ���;������~�ޑ��+�.�=̞|2�>;�������6"""""""{kQ� DG��ܹ�j�4�=���R�۟3�>��y�ڭqmm���=�;f�X����a�q�S=Bq�r:t��*�quuA\\T���<�=:u
�'��ސa6�@ �GM���0}�W8u*�nc!""""""��zt�\c1S���e����h���2� /�4[����l''!>���ݻ5�N�.��m,DDDDDDD���B����R\�P}]�a�:C�����+u�c��N��5|���ô
��	_}�(�wÔ)��n��5�z��������z���!66�^K\^ye�m;W�N1���Y��+CTT &M�		YvQciq� t�R�0���k��:��޽#�x��Ѫ�Rg�^�$""|1q�2$%��{HDDDDDDD6�"C��]�_}1S >�3rr�q�Db��y��{w<N�L����$�9����&|�[���=$"""""""�j��G�.!�j��|��>��
�����O�>������^�[�\.��uO��C����ɹ��ʹ�УU+��Kj��eǎ���0{�8|8�]�w֤PȰ~�lxz�b̘��~�5>�������1����T�4��U_�0m]���S�6��    IDAT���t���C;a�"���0��t���� ,���-�q�^""""""��E� �C��gzDG� 0У�K\ Sm�S���{w|�۰6�R�Yh�>���ӧo�{HDDDDDDDV�bC���P�ǧA�7T{�@ ���ض�\����1�Fu����`4�}'[��L���Ɔc��e8v솽�DDDDDDDd5-6���%M��L`��n�p!7nd׻��^�K�Ұ}{�g�؂D"�ʕ���v�:�8p��C"""""""��zDF�������\ףG�y`˖���M?����[��K�X�/������W`׮�n%""""""j*Zl�!
Э[8N�H��X�@�솭[�4��W_���|�ݡ�cNNB|��TL���?�V�>l�!5H�= �W�V8u*�Vǎ��/��ʕ�z���3���R��w;���$ĢE���c����5�$DDDDDDDuѢC���p\��	����c�uEX�w�g{̞=�K��lP;�4o�0|��,_��?�:]���DDDDDDDTg->�0Q���%.�� R�3���o�9����F���{���Ν���#_�*"""""""jJZt���!Cd�/N�H���GwCBB.^LmP�?�N����[[Ԏ��͛�ǵkY;����{HDDDDDDD�֢C �ٳU�C�.]Bж�?6m:ՠ>,x;w^����Ԗ�u��_����Q�>F||�[�5=zF�̙d�+�9n\,~��d���J�^�5�+,���l-8��7�AD�7F����uM�������C�=bb"�T��ڵ�Z?n\,���8|�Z��~��Q�z56op[��P����1aB̚�o��ee{��������J->�h��r�Ǐ'����P/���
?�|��}��y�'��~CI����ٚX�����X�d2��� �M���%�Q�Z|�!
гg�Z� ���=��og�Vk��ܹCQVf�g��ip[�eҤ^ز�y\����'O&�{HDDDDDDDwi� ���G�&����
���v]lp��������}HM�op{�%::;w��[�b��O�ᇻ�܅�������� z��DJJ^�C�B�!C:��OX���S� 2�l�J{������,�O>���}���<{������� C @�na�H�8v�F�ϙ0�'�ￂ������$�{�Ƕm�w���ט{�?�m{�ť����EaV""""""r|=`*�^�%.C�t�\.��l���L��o����*m6��mۋ�<�7��[�iӾlV�u��������0�(קO�:������ñ��cV�o�BA�
�}��jm6&.���Crr.Z�o�9��X�9:]ΞMi�QQK�У\�ޑ�v-�N�U&M�+W2p��M��������H,]���s�Ҧ=���?�x�=����&��)�*=v�ܵx��%����{5=���F@,v±c�_�ҡC �u��l�)S��s�`��_?Y�M{pq��Fb���Vk1x�b��ί()�X���)�Ν� ��+֬9b���b�QN*uFtt(��� �4��l9��R�U�!
��{��W�i�)��iO�:���a��1���0�=l�r ��'�C�7msk4����/g�9\""""""r =nӧO�:3�1c�C�-�o����8:u
��OonB^^��ڵ�H��3������g���G�o�=���r��<��wط�y�`CDDDDDDMC�������iu

x�~��/�������,\�Ū�ړ��+�,��-[�"3�����F�F��>�5N�L�� �������a0��M�^� 9�Сku:oʔ�8t�U��J$b,^<?�t��_�Z�M���iiyfy�F��L�����v9
���J�^����{�""��o�B����ŤI���k�Ri�ڶ=-Z�Ba�?z����}����F9�w�ׯ-�[�!����?�t�BC���h�TZ���oVm�^.\Hů�������PR���qK��^�H�#""""""G������Í�HK�ۅ�ĉ=QTT�m��Yu<2���x�\�'��[�զ�?. �b'��N��ח!7�&|�����9��h4�{M�NW��_�;�<��{�����������>�g��g���￿WW���X�J5�����l$&f���t$$� '��i֌X섲2����<=]q���˥�:53=*1mڗ��r�'�<R�����Ǝ�����6m��:��|#Gv�;�<lն��J���l��3�D"O���
= : ��((�f߁6a����h4�Q��У˖�Ŋp���|�A�0`@.c�q��u3g�ď?�B�~��~S 0f�L�:��\I��٥����Ml��5]k׮��͛����������&�� ���᭷~���Yu��1}z_,^��珄Db��a�:c��x��������.�j�Mń	0a�{�Y��tؼy���ADDDDDԤ��i%:t����R�s~���2l�r�#���1�j�x���m�>��`�Q	�P���o��:�+�K1qbO|���P(d�䓩ظ�͂"""""""G�У
�w��Cס���|�����4>|�#��k�Y���W7�֭|��ADDDDDD��1��Q�ht8r$���k���(|��A����WG ,�s箩��+�0������t	���u_� �?> ;v�Gj�mfb��N����8s&�}��&}4��^�5�X""""""jzTc��س�~�ǠA�⅕+����֦��|s4���8~<�f�5G=���W3�5[C(��'���Bi���3�1�^�	�<���Kl�Qs�У���˥��� &N��F��>a�U�d��DB<���F����U�LE �����QS�uy�����!"""""��1�����qqQس'�^绹�`��>��6#�r	���Q8p�������l~�h4V�z��}��f]^k�x�������j=j0p`����^�?�Tn����_���*��%�������_7l�WSTY��VaSC��ν����h�3t������l��G��b��_�쉇������;�J̜�#FDc֬���-�yMEcΌ0�Ĩ�R���GDDDDDD��У��rt���;/Ի�����Gp�d�GV��ߟ��O>�m�g�47��,��e*U�sy�C�Z:�v�T��;w����|�^+��r��|��c�p��z�����Ե�GC� """""��c�QÆuFRR�����ƬY�}�9$%�Xqd�k�. }4_�'֯?n�����
��ow�ب�r�;ϫ�ͪ^�L"""""���У:tDX�7�����H�BǎAX����= `Ĉh̝;����s�R�O{�3@�3h�nIIM�W�gmڬ���Y�{""""""��a�QKC�vjP] �={06l8����)2��ޏ{�i����E6%""""""z�ڰa�p���>�
|��>��NNB|��t��Nx��-��iCܾ<��5/=j�O��pss��]���!	1g�|��A��8�����]�4�]�ļy�t�w.y�+DDDDDD�C�Z��0p`��G�wq���{��C���>`���,"�+V<��[�`ɒ]��/�=1�����;c߾�P���nC,v�3��W_�RYj��U�_��x���X�d'6n<�h��C�:2�##��oP;S��T�o�=h����ԩ}�쳃1o�:�:�ܨ}56�u��.������gԎ���<3_~�%%+��v���A�:`ƌ�~=�Q�&""""""jL#+4�������?������"�w;j��{��ٳc��AVa���4i9RS���s�Ѩ�WǼKʄ	�<��eÆ ���DDDDDD��L�:>�34=��m���O?=˗�JU�!������Ӧ}٨�Ej2�|�0a�̟?��� """""jR8ӣ�M�^^���GԎJ�E�>o��'�0g�}V]�`Ԩ����gC*un�1�
gz�èQ]�k�h���#�9�������B�T[it�h
;��r0{�w(+34��������l��G=�g��:����m��}���e��Zadu׺�V�z�y�=�=�""""""r=����}����m�ܖ����Ê��Sl���]LL8V�~�v]�?���x""""""�握G=��;v\�NW��&M�__w|��VY��{o|��Ll�|������Q��У�F���J����H��_~ �VBzz�FW?�Ǌ3�a�q���FDDDDDDԬ1��'//W��EaӦ�Vi��U+_,Y��*���}�uĲe����G�p�DDDDDD�l1�h��cc�s��T��%
��k#���p�j�FW#FDc��iX��O̟��""""""j�z4���w ��y�*����x��Vi�!F����u�a�ܵ�Յ�������� �9���;[m� ��?a��x<x�jm����w���O���a���V)�JDDDDDD�Xz4�ر�ؿ�
��J��^�nax����i[���Ea͚���<��J����=$""""""�Za��@qqQpw�`��3Vk�_��k�2��O'��fC���?�0'N$�G�@A���C"""""""�C������ݰi�)�����E��A�nx�Tk��=?��n���ȑ!11��cY����������V0vl�Oĭ[�Vk���B����/�[�͆��!��6^^�9�#9�p�1Z����D�~�����C+�ٳ��=�y��f{������������(�Z���㆟~zqqQ�<y�/�WaKە+ n���o�l�a�i���=��N  ?_�͛Oa��~Vk�s�l�x�/�c�ȮVk��D"!F������m�ɓɈ���Z��c�}m���ܹ[pq�W�H;��������Z"�����ޒ�sѷ�;زez�he�v���?�ƍϡw��<��g�Y��]��`Ϟ������V `��G0n\�GIDDDDDD-C+?�3�j��ߟh�v�~z�_��Ν/A$jz+��J5�y�;��w��mv@(⧟�m��9��w݌M��[���Je�W�|s4��r�j�A��k-r�%%���^3M�G]���;��������Z*�V4rd4~��U��ļy����;��[lն�aǎ����*wk1()�bϛ���������11��"��=����z�O=oo7���/Vo�!�Z=���M�=ɣ����J<��P��;��������2=�lҤ�8v�՗r8;��p�l�p'N$Z��8q"	��� LEK��ח�ҥ4̙�,%CDDDDDD��-k�,(�[��Ai�����jۑ���t)6��ԩ}��d��* @�v����D�R��R @,v�@ �pF$$dA�ѣ�~�������n��[l`ٲ�X�� ������^��a��Ax�aVm�Z�����Rq�|*ΟOArr�ʌ
�^���'���h[�>}� 44��� """""j=l ;�=z,�7�<���;X��o�=�6c��Ѻ���۷�F��Sgcǎ#�|���*�9���Z��3gb�ʕ�Q�`�a#O?�
Z��|���6�3f)��ظ�ki4�<� `͚5vI���?�4�/
ᠦO��w_���&�P�>��S���f�Q��ODDDDDD�z�H߾��g�P�]� ̙s�~{+23m�Qs���F�Ok�@�+�I�?���x���6i��������9c�aC���@I�۷��I���"���D��q[���IDDDDDDD�C�˥3&�V�Y�zE�'��~BF���1���3�ő#	�z5�f}̟?
��r����f<DDDDDDD&=l�s�`�Ɔcժ�6���E��K��Cװz���!""""""jNz4�3�᧟���Dc�>�t	�/�[o�����������~e��|���j�m�f��i���P���D=��v�X��˦�̙s�����kQVf�i_�I �h4�h4Z.�o\�qw�V����fM�U�މ������n=���ӧߋ+�`�]��H�O>y.����Y?���:%��[b���k���j�5[������j��G#�1�^������/ڴ�֭������;p��M���(n�Ab��-5�Y���GDDDDDD1�h$��r�����o�{�?l�Y�VA�Tۼ?GPݒ��_��Lk,�!"""""��c�шf��#Gp�l�M���)��x�mڗ#�ˌ���m�3=��������G#j�>qqQX����6<=]�l�?�}�y|��!���ܹ���ZU-��y��}Q�6�,�JDDDDDD��У�=�T�m;���|��իW$^zi8.܌�Smޟ-�TĴ��U-�n�Jmϫ�������WW䔡Q�z4���(DF�a��?����^�"1k�j��h�O""""""����G#x��X��h��NNB,]:J����d��Z�ۗ��y#"""""�����<�p�DB�]{�Q���s�ҥ�`ӦS�6���ݹT�;�5==�@"���cٲ���������+`��-8z4�Q�$""""""�'�v��PR���u�������������/�=0���\�3��������=�ʲ��o�kP�R2��XF��v*Oj^r����[
4R�@-!��a:���B`�m���%B3GH	oa�0.��%ܗ����!׽6{�w]>��5{ּ�}��r3���<��FssKN�L�Rq�-�ⓟ�+��9�   ���H���'��o��g?��9;w��ɓ/��^{'F���ټ   �kJ�u���8����n�--�; �G��1i����:�  ����Hؐ!'�ʕk��^��'�����3b̘�b��Ws2guuu�����q�^����������  �A*����ꪺx���1w��J�r6o&��a�fƼyKc���ѳg��o��ձhQn�ˎ{�q��'   '�y`�ʵq�	�bʔ�ѫ�s:wSS:���;�/;{ldp@���   ���<н���o'���ܕ��q�����"�76�<   t�G�>�W��ª�?���Ͻ����Kb�ʵ1d��H�s�]   �HJ�<��}�7��h$��G��1mڠX�������|~   hoJ�<r���/��f<�ȒD�?���q�ČO���O$   ��G�ѣk|�;_������l1����;�O\��1k�'�   P��yfĈޱfͺx��g�0`�qq���G?���~!�   �'�y�����.:!n��w��؜X�+�8-�F63�xbib9   ���yh��S��6�̙O'��'?�f�w�Wc��_��&�   ����C����<����'��hL,G*������8�/ǀ��sϭL,   dK鑧>1�閘<��Ds����ĉ����|��W,]�z�y   ���yj��>�^�q����k?H4KEEY��ߋ#���;Ɋ   
��#�]t�	��ޝ⦛~�t���,�i��׾�/ѷ�X���~n��Q_�|��  ���y���"�����1��x��7����q�=��9�?�1gΒ�\߰�!�>��:tz����$�   6Qz乳�:"�:�{��P�Q"b�V�[o��\2-n���Ғ���	����H�W��?o   �Ie2�L�!ص?�iU�y�-1}��q�)=���ŬY�b������.�}�����N��e��>�b��+�[�}N
  @)Rz���gƻ-��  �IDAT�%�c��EEE�,�y1h���ԩ*֬Y��-[�UT�GϞF}���ԩ*��   �����]=��X�f]L�����|�1�t���W�\��G
�����t��/oĕW�:�t   �2�G���m�:��?��X�~c�q�X�nC�p�c���B�tK��?�&�>��   (yJ�2t�)Q]]&<�t�-ƍ�64D��wIe2�7nN̟�R�  P��S��=�̘:ua��J�}���1s��������X����
   6Qz�s���8��CbԨ"�3h�t����~ѹ�CJ��RQQQ��϶�d��!������˘   �(Oo)@/��F�v�Mq��E߾_M:N��dbٲ��V�/��E�V���oE:�����H�3�Ҳi5HyyYwܡ1s�%Q^�s  ��(=
�ر����/�'������l���8�-[�t*6l����+����b���hj��*���n�/}����C=4ƍ�t  �v��(P64�I'�'�xX��7�8[�R��������ZccY��~u��V�8�������ShJ]]]]DD�[�   ړң�͝�?q�S��~X|�+�M:NDl*=fΜ���K:
Y�������+=  ���P�ֻ��q���F�ESS:�8   �W��g?��V�o����t   �+J�w�A��ȑ�c�c͚uI�  ����(��ݻw���~g2   ��Sz�����0���?���������O{)E���  rA�Q$�8���^1f�C���ʔ�)K   ZG�QDF���_\~�}�   J�ң�TV��ĉ��\���T�qZe�U�Tj�+�1��og��l�ּ�v���om�m���   �J�Qd?��>�W��H�Z�6�8YI�R��d���->��o��{:Ǯ�k�ܻ�y��+y�d~  �b��(BÇ�=zt��#g�6�l�o�َ���5���ٺ��\j   ��G��,�[o��>�ט2eA�qZm�U��ZawْΝ��   �H�Q�z��#G���4V�x;�8����4v�m�kI��Hz~  �|��(b�]�+;��2��hjJ'g����Z[V�S�˕lK�|��  �KJ�"VQQw���X����ON:�nm���#V,�j�]ma��lr��}�1?  @1Sz�C�?n��<yA<��Ҥ�lgG�f�Ecw��f3Ǯ�����lr��}{:?  @�Sz��o~�����1bV��ƻI�  ��Pz��1cΎO}j�����N�$'+[o������$��*   {N�Q":u����K����o��t��l��P�r�I�B�~   �N�QB;�����o�ĉO�SO-K:   t(�G�������).�tF�]�A�q   ��(=J���}���<��^p�{   @k)=JP�.�b�ԁ��s��{8�8   �!*�@2���O��7;���~P��|��Ʈ������v��WWW�t  �v��xDDI;���2eA̞=,�8��=���:�!�VUUI�   h7J��N���2^~�͘;����O$	   څ3=J\yyY�u�w���"�MM�#  @�Pz]�t�)S.��K_�����I�  �v�� ""���nq�-�bڴ�b֬EI�  �=��`�3��r�qj��@,\�j�q   `�8Ȕ��d21l�̘7oi̞=<z��t$   h��ijJG��w���oǜ9?�n��I:   dM���_�a�sέ1{�����c	'  ��8Ӄ���c1c��x�ݍ1h���  ��(=ةn���3ǋ/��#j#�nI:   ��҃]�ٳ[�s�E1gΒ���$   ZM��n���替���T�vۼ��   @�T$��Ч�1�v�q�EEEyr�?������Y  �<+=h��/>1����;���4���]�1����g�翔@:   �(��%kS�.�k��#F�W^yZ�R�x�����_6|�;WǼyWF�]��
  @	�҃�]x�	1~�yq���c������W_�`444FDDccs|�{��ƍ�	'  ��Y�A�-\�J\|�����|��?r���,�:머��J  @��҃6;��������__ee��\knn����c��'J  @�Sz�G�oq47���e�C�L&����X�xE�   (uJ���g_�i�Fss�.?7p��x��9J   �(=h���t��{g�R��\:���a85��ҹ	   �������wc�Ʀhi�DUUyD��hnNǒ%����]@   J����f���<�Z<�̊X������DSS:*+�#�n�T*��~~�s��	%  ��(=h7��ͱd��X�xE<���X�xE|�AC��oZP�No:���GG�QG�dT   J�҃�TWWGccc+?�������꠨��tTWee�#�i�7߼�Cs��������!�   ��� +�T*�>���ׯ_��_��!��SѥKU;'�#���F}}}��  PH*�@ᩩ������c�CMMMQ__�t  ��xz   P��   @QRz    EI�   %��@*�J:  @�QzС����N  �R��    ��҃�yE��?������Tj�kG������d;���w��5��&K6�u��  ���P�2�L�R��d2Yݷ�=[��յ�s��n�nَۚ�/�q2�L�'   ��Jrf����#|��m��Y���]��eB6�e3  @��҃��uQ��}!j��%��   �҃�Ӗ�-���2�w  ��[ȩmϔ����|_!іq��;  *+=�pٮ�����no�1w7���i���d�B]!  ��jGX��Ύ8,�-c�.kk���p�l�k�8�  �T��   %+=(
�:���  �Ҥ��(�C��   �'�[   ����    ���   (JJ   �(�2N_$���RSS�pr���."�
  Oo!+�G��e˖%�����C=4�   Y��   (J��    ���   (JJ   �()=   �����/g]��    IEND�B`�