�PNG

   IHDR  �   %   ȥm   bKGD � � �����  �IDATx���ALW����`cՃҤ۬�&�i�z�5�&���EC9J���H��p�Wbz�`�f�a�]���h�h��
Z�Zl����
���Kv-���3ofx��ߥ�μ�}oƝog�몬������H^G�΀���*3""��I�Ō����վ1;;��Ǐ#���	v��a��׻��)8���i��񠫫���n�b�ɓ'155�vB��~�>}z���v5cOO���QSS�Tnd���a455!���)����������N�򜪪hjjr;SE �?K�� t�]sg�t��)S"'x<�S�L�bL�#Yd&s1NJ�l��I�Ō����bFDD�c1#""鱘�R[[�h'��;+��0�o�c5#��C�q���R�x�Nmhh��R�Fc��Ǒ#݈D�q;��7��2z<�@�������C�ի?�����<w)��S~����	��'��  ��a��w\ΎH�?E(4U�ѣ?  ��O�w��.g�����Z�y���.d�6�w'z}$_kcj�L/]�ڶF�4O�_��H$V��Ph��(���[�����՗�7{�o����'�+��ھ��z�k�Zݖnz9i��&^�>�mE�O{��!�Zo�l�e;���00p��=&&f�����I[����L���߹L��*awfz�Fo��k�1��3ӧ���1�T&'g�AUØ�[���yU�r��i?xz��^�W/��mV��!j��Ɨ.�^?z_"R��&7��aq1���	�����[S((P���=W>G��g��M��*a�,������ؑ[���۲�W�Hă���P�0���Da���2��)`���hd�LRm�9�`��l��S�-�}E�� ��x111�k׾�����' �|ʑH�7�g��si��13rr�L��SD����L�.�y��ܻ��o�z/Y�2ih��Rl6mڌ]���i��T�j���v�szv�:��ң��~�u�˗�"˺�h7~hk��a�iN3 �<�z��h<36lx��������̃X���X{�g���Y�o�ٳg��iׅ����G+N�szv�2����PYل'O"��P�D"c��ʷ�����|E:p�۶���i:ɕbfw!����nn�O*(���b	��Wx��w�Bc��cv���7ꩮ���j����V�yĨm�n��~;�:.V���j�h������������x�n����G���.+{����+���#qܼC�������}D�mgT�x��4���L��SOEE::>ǉu�F(4�K�F��ً���ֻt�dV5�kkv[6���S���i�ꭎ��K��4[�JJ���X���*��?���]���16���x<	oZ-ўG��̌,x0{1N�.SL3�.2�(�Om�2�,EQPU�CU����q�!��Q\�2�H$E���fd��կQF'�E�)G}�*Nٶ�㸘�eK	ZZ���R��������7��g_�^Z�
��l���N�?뽶�?g��<���T�̙fLN~�s�Ğ=� ��7���<��7������H�� �c���2��\] ��q�z�٧\T\�E]�N���t;����Q���+�۷oC{�>���s;���j1c��|��+��O��1#I�Ō����bFDD�c1#""�\ 2<<�`d���:t��4,QUn�A$=UUQXX�v����rۚb��� ����eD���|n�`���C,�� SnH^eTTT�P(�P(�v*�龯�p�,��(�̈�Hz,fDD$=3""��I�_�eD�l�    IEND�B`�