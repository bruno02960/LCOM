<map id="read_reg" name="read_reg">
<area shape="rect" id="node2" href="$group__rtc.html#gab7e8ff751e63b72d14aa5f7ec727d337" title="Returns the day on the Real&#45;Time Clock. " alt="" coords="132,5,195,32"/>
<area shape="rect" id="node8" href="$group__rtc.html#gad751c36263a847ec77044899618cfd66" title="Returns the month on the Real&#45;Time Clock. " alt="" coords="125,56,201,83"/>
<area shape="rect" id="node9" href="$group__rtc.html#ga37f344d06f4e1b826aed5adf7b729fe8" title="Returns the year on the Real&#45;Time Clock. " alt="" coords="130,107,197,133"/>
<area shape="rect" id="node10" href="$group__rtc.html#ga57e0eac5ae1c791f2c63b0740ab94e08" title="Returns the seconds on the Real&#45;Time Clock. " alt="" coords="132,157,195,184"/>
<area shape="rect" id="node11" href="$group__rtc.html#ga59e635249f9555c53ddc24e54b82f01f" title="Returns the minutes on the Real&#45;Time Clock. " alt="" coords="133,208,194,235"/>
<area shape="rect" id="node12" href="$group__rtc.html#gaa14f12da2be63f2a594cadff28d10f40" title="Returns the hour on the Real&#45;Time Clock. " alt="" coords="130,259,197,285"/>
<area shape="rect" id="node3" href="$group__file__handler.html#ga90d3bc0149cb0d2782d63aa42cf3fa86" title="write_score" alt="" coords="249,132,337,159"/>
<area shape="rect" id="node4" href="$group__game.html#ga02fd73d861ef2e4aabb38c0c9ff82947" title="Makes game initialization. " alt="" coords="385,132,424,159"/>
<area shape="rect" id="node5" href="$group__print.html#ga92978930f74831bae9a6d6f22d089615" title="print_menu_kbd_or_mouse" alt="" coords="472,132,651,159"/>
<area shape="rect" id="node6" href="$group__print.html#gae91d4cbee2dab64187187499dd0eecd4" title="print_menu" alt="" coords="699,132,785,159"/>
<area shape="rect" id="node7" href="$group__spaceinvaders.html#ga3c04138a5bfe5d72780bb7e82a18e627" title="main" alt="" coords="833,132,884,159"/>
</map>
