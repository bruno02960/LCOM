284e5074e8066b7270425b43a1f9c232