<map id="object_creator" name="object_creator">
<area shape="rect" id="node2" href="$group__game.html#ga02fd73d861ef2e4aabb38c0c9ff82947" title="Makes game initialization. " alt="" coords="468,34,507,60"/>
<area shape="rect" id="node6" href="$group__game.html#ga1fd9e64dab3abe9facfb4dd7e1267bae" title="Creates the pong and switches game state. " alt="" coords="184,34,259,60"/>
<area shape="rect" id="node7" href="$group__game.html#ga671b58f5509a3a9fa692bacccfc32cc9" title="Receives drivers interruptions. " alt="" coords="333,84,420,111"/>
<area shape="rect" id="node8" href="$group__game.html#gaff72f275b5af37960b3baee51f855041" title="Makes a game round, where updating action on screen. " alt="" coords="194,135,249,162"/>
<area shape="rect" id="node9" href="$group__game.html#ga425ea598437d36368c0e136f2be75a61" title="Makes enemies down movement. " alt="" coords="157,186,285,212"/>
<area shape="rect" id="node3" href="$group__print.html#ga92978930f74831bae9a6d6f22d089615" title="print_menu_kbd_or_mouse" alt="" coords="555,34,733,60"/>
<area shape="rect" id="node4" href="$group__print.html#gae91d4cbee2dab64187187499dd0eecd4" title="print_menu" alt="" coords="781,34,868,60"/>
<area shape="rect" id="node5" href="$group__spaceinvaders.html#ga3c04138a5bfe5d72780bb7e82a18e627" title="main" alt="" coords="916,34,967,60"/>
</map>
