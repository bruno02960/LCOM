�PNG

   IHDR  �   �   �{��   bKGD � � �����  �IDATx���{PW��o���@LD]|� �|�Q1��a��M�V����Jv�*���w���ucU����Q#�Y^��/�K�eU�#@ķ`d������0O�g�������>�s��s��iAEDDD$)��2�,0!� 2������߯~�+466J��mܸIIIR�A�˚��M �V��8����Gvv6����$�2���<dggK�l���HI�א���d�	���H�����d�	���Hة���V_�nS��\�W�(��M�jL�D�5A�,�%Os�U���9�M�DDD2��LD�$B�i�sߴ��[�ז��{?�_se����8��dMD�c�Tli���}�xM���%F[��M˳�|=�{"[0!���L���ܝ0���L�D�q��,�Ȼ0!�ǑCT1�wa�."���j�r���!�|�!���10�{?��V�ʷT��񙋁�L�D$K֒��i�
�hy����L�b�5������LD��&a�EL�D$KL��k�dMDD$L�DDD2��LDD$L�DDD2�N]D䔎�n�����w�v����������P|��!��j)B�����j�R�AbB&"�]�ֆ������BB��� dem������y��S�JI�	��l�o�2}CY��Zlڴ�Qy^C&"���?��Ji��*��ƍ#�aӦ%n��ȳ1!�]23�`0�9�R�������@t��a��ȳ1!�]f�Cp���(�����O�	��)2"��k�D4��n����QVր#��V+��?\S������W��";"�%"��CAA��k��މ����̌�̙���Ǉ�U�P��رc�$���s��LD�v�5��N���:f��+�$ ==&<�?_dd���(B�����""�0z"��2��K���z�t�PQq��#���6��M1�Lnn9�n- `��aϞ1nܨ��ȋ0!�(QQUu:�)��֣�K���h�<��l��Yo@�s�>"#����FcǎMP�m����cB&�1�/�D~~5������7=ii1HM�AH�}5���`�H�!�����|@{{�Caa-��."44))��k�D2��L�zz�����(,�Aii= ��#���+fA��0DrL�eΝkEAA

jp�Zbb������:<"��	��ܽہ��Z�tը�oBX�ddh��j"uxDd&d"������T���~~*�[7Z��M�B�Q��<	2����o�NW���:ܹs��3��j�f��x&�`L�D�o����Z44\Ō�HK�Ezz,���H� 2�Luu�q����ĉs

@r�<h��ĄK�2�����S�.���%%u�����'GFF��=��<2�45�FAA��q��MDD<��̅X���ѳ��3��6�D����>;����.bܸ�X�>��9z�b�h�"**.�?��h���V���g�D>�	�h46^�Nw
�ŵ������	�V�Ar�<�(uxD$l�&r���N�ުT[{aac����tf��:<"��DUU��/_[�n5�
=�֭[%�����V���>��8z�3���|j�"����'��'�WUUՠ�mP��� ��_��t�x뭷p��%��pإK��V����'u(^���?��-����������n��� ;;[�Pd)##������{�s�M�+V�pwL���\����j��j���8x��!9����DDD2��LDD$L�DDD2��LDD$.�y�ʕ�?~�UŒ��qf�M#"rK癁��`vY9��\RC^�r%�?����u��=L��*�{n'JK����A�q��n�@����!r�O?��ĉ��7�PSsIIk G�AQ��p<s�./p�� ��'���/�c�5֮�Fjj�-{J%�L����� ��+�k�I<��#��� %e�x�@q5���}Mզ�Z�����:�-g�L[�3��S����::�q�`��?Ĝ9o��׭ �/k�M?��s�����W��u�+�U�سN"�*����n��mر�8���e����;����.[�=Ǖ��){�	��t�����M���f:���l-g�2mY���)�� p�n�C�n���_��>�������\�j���}MJ���p&NG��=�'�;�\�x۶��o�":z2��X$%����Av�i����W$IG��r{����);Z�-����pĭ[�8t���u���;V��u�s�q���1�����;ӧ�si,�N8�*ϴ[�u��Ǒ�nޔ~�"���p�v[Q���\_߄�g���ň����#�;�Ng��Z�X{oi9G��a���m������K{��f}�n/_�	  ��wI�ܚn��#e�������:M����71}�M�������bp�1hK�Zo��<:!{[/�ŋoJ�p����X��!�S����{���X���aĈ�a�p0�5��z��p'�eˤ߿�w}�����w�X�G �R��N�V�V�����p���Rӷ�uzl��5�^CvG�J�R�`����AHO����1�� ���8�^�q��3ן~ND��j�z#"#à�j��<&< ��~�p�CgR�Ű�o�+kB6�VkO�����-Ӵ<oJ�*���� ��.@jj4��P(�O(C5��Ҕc�[ʷ�`��Y��x�]��;�������m�����8]����U�[�o˱,�&k�i�ok�9�G>�7Pc͚h��.��峠V+]�k���2\U�������Y'�܉�����N��Z�\�.{����<�qkOYCMs����&��6m�x$'�Ú5�X�:#F�Iy����?6,vY+�9�%��,���bw%Mg�����_��;��:�6C��\sx`�Fdd�?�����^�H�C%Cw&er/wX�z�y+�|�"�,0!� 2�0!ɀ�N]���o�3�t��	dggK�S����^/u^Iܺ��c��P��a%??���/�ݸw�mm��w������O~��;?�� ��u$fϾ��@�ԡ�ڠ�������,��H3Ʊ'�j���ʒ:�eee1�ѽ{j�;7J�!!��0�AA�6/���y�ݻ˱k�I�TJ���&���n?Hb�����Z���j&����BBB ��}͉��ڵv|�it�*44\Exx�Z224#uxDvY�������+A������#�L�D��̙f֠���o�ǢEӡ�j�n�\��/uxDC*+k���`贡T*�R)��G/ !!���y&d�a��������58z�,�j%�}6�鱈����	��e4�X��whi�cu>�J�#���'/a��St��	�HBw�v���������+���X���bƌP��#���a۶Ã��Q�		B~�˘>���=���d���:t�S(,�Akkbb��AR�<�(ux��.^��={*��}���ل�R)1uj���1aB�Qz6&d"�1ETT\�Nw
���0E$&F!##˗ςJ��hx�"�;�ݻ+���0y�XlڴWQRR���w�(�J��L�޽����F���d��/9����.bܸ�X�>����ᑗ�}�>�=hi��'���-[�bժ�P(���-X�z[��
��g���?�i#��e��"�ĄL�!�\����Z��W��囈�����8�_���QR�G^���&��]������YYqx��xL�:~мk�nG]�w�6-������7�`B&�0�(���"
kq�P:;�X��	���"11
~~����()���'QW�""&��"55��~�+)��O����3x��a��{1!y��.=JK�QTT�/�8��� ���GZZ,bb¥�d���������
��X�&[�,��lZ^E\�چ�G�9R���L�%�]kCAA

jp�\+f�EFFRSpT0ЛD+*. 7�G��EH�(lذ6,f�h`B&�B��M��Q\\���N���Dff�8*��w����-Gc�u,Z4�7/Ś5s�V+����	�ȋ��
v�@����ºus�����A8*�7;����(,���("--�7�#"b�ԡ�L�D>�֭PRR����M���Z��C��\�`0�=�ݻ�QQшi�����㑙���R�GV0!�����(*�EAA�_oGll8�Z����u����s�����cG�1Z�ō���W��?�ĵkmx�Hl����g�%�C0!���#N�8���>| ����tV��e�����*ށJ��ѣ?�Op�)��\Bnn9>��4F�
�s�-ĦMK0e�8�C#;1! ���%%u((�Au�%��#--ii�fG���J��' 
��)�s��x��H	"�=]]z�b��
�9ӌ�s'c��HIY���<2r��M��W���MM�=��$%�GH�(F̛�&n߾ �M�[����/'H�W�r����'�T���II�e�R>��K0!�E}���t���g���m@BBf����Ga��zA��� ﾛ��\�hq��?�{w9����c��q���,¸q2՛0!�M:;�q���t���7M��|`�|J�QQ��g�O$A�ޡ���=�r���gb˖�X�:�cF{)&d"�K{{���
��������}�^BTT�0F��ΞmAnn9����J�@z�[�,Ō�R�FnƄLDvٷ���^ ��rBzk�*�|�k����<�^߃��z��u�՗���b��HO�ŨQY�W0!�]�}v;N�n�-��B�(?�y"^}u5�5��چ}�*�o��p��}�^�-[�aɒ���|2٬��4��:����o��D��Ѵ��kD}�-��x���O��ѽ�a�R���d�T��1������R�![��/2�L����~�����cQ{{'��  Q���  47�������B����� ���/3��+��_EW��bϠ����HII� 2��G���m_���ED�P��رc�M����  ��r|��QyA���!uN���Cvv��aȒ��˾�DDD2��LDD$L�DDD2��LDD$��ED^O��&�5�6�n���֐��Ȭ��;8�U�0,r��*Q��p�k�DDd֋/�3͘>=Z�))�1e�8��2�/����zJ	k�D$}����A�_��j�#�7�~`l��3��Hr2v�H �ŋױm�,^�َ֬]�N�ƍ{.]������k�57���w�sk�D$+k3�5G��s�X�2W��g�}噛�S��������7���f��f1/��V�g����� ��ci{Y���m#s�9��;��9�	��d�֓�=�&cm���<1�BE�����oQYو_�R�U�f#==�V�v�|w�*�+������̄LD�f�����k��E����/��#Y p��]}��4{������#g  �<�K�pe+G�<˶t��Z���r2ɚ����CW�dN���g�s;X�ֶ���ɚ�|�����Z������ƍ�%8Cv��hi�kq�B�  B�T<�d��C�j[ڲ\����5dWbB&"ٲ�<8p���I�O��:���KA�R)�h�x�t�t�g[Z�h���M���u�ɚ�|�P���MsE�*[ʰ�3o����Z!�T*��cDt�dh��HJ����\�.{��rG��]�	���̺}�> `�4���������gXk�fB죏^@k�]��Nu�z���I����g8s���$1i�L�4fX��߯)�IDD$L�DDD2��LDD$L�DDD2��LDD$L�D����ؿ�Cώ�˶ J�����#��(�`~�
"���455᫯��:��T*�����3�L���Dss��aȖ��˄LDD$l�&""�&d"""`B&""��פ������?>�3�Ѳl�    IEND�B`�